-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    num_cont : in  std_logic_vector(15 downto 0);
    row1 : in  std_logic_vector(15 downto 0);
    col1 : in  std_logic_vector(15 downto 0);
    rk1 : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 96)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal num_cont_buffer :  std_logic_vector(15 downto 0);
  signal num_cont_update_enable: Boolean;
  signal row1_buffer :  std_logic_vector(15 downto 0);
  signal row1_update_enable: Boolean;
  signal col1_buffer :  std_logic_vector(15 downto 0);
  signal col1_update_enable: Boolean;
  signal rk1_buffer :  std_logic_vector(15 downto 0);
  signal rk1_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_46_branch_req_0 : boolean;
  signal phi_stmt_48_req_0 : boolean;
  signal phi_stmt_48_req_1 : boolean;
  signal phi_stmt_48_ack_0 : boolean;
  signal n_address_282_50_buf_req_0 : boolean;
  signal n_address_282_50_buf_ack_0 : boolean;
  signal n_address_282_50_buf_req_1 : boolean;
  signal n_address_282_50_buf_ack_1 : boolean;
  signal phi_stmt_53_req_1 : boolean;
  signal phi_stmt_53_req_0 : boolean;
  signal phi_stmt_53_ack_0 : boolean;
  signal n_word_start_271_58_buf_req_0 : boolean;
  signal n_word_start_271_58_buf_ack_0 : boolean;
  signal n_word_start_271_58_buf_req_1 : boolean;
  signal n_word_start_271_58_buf_ack_1 : boolean;
  signal n_winr_211_72_buf_req_0 : boolean;
  signal n_winr_211_72_buf_ack_0 : boolean;
  signal phi_stmt_59_req_0 : boolean;
  signal phi_stmt_59_req_1 : boolean;
  signal phi_stmt_59_ack_0 : boolean;
  signal n_left_290_61_buf_req_0 : boolean;
  signal n_left_290_61_buf_ack_0 : boolean;
  signal n_left_290_61_buf_req_1 : boolean;
  signal n_left_290_61_buf_ack_1 : boolean;
  signal nl_start_37_62_buf_req_0 : boolean;
  signal nl_start_37_62_buf_ack_0 : boolean;
  signal nl_start_37_62_buf_req_1 : boolean;
  signal nl_start_37_62_buf_ack_1 : boolean;
  signal phi_stmt_63_req_1 : boolean;
  signal phi_stmt_63_req_0 : boolean;
  signal phi_stmt_63_ack_0 : boolean;
  signal type_cast_66_inst_req_0 : boolean;
  signal type_cast_66_inst_ack_0 : boolean;
  signal type_cast_66_inst_req_1 : boolean;
  signal type_cast_66_inst_ack_1 : boolean;
  signal n_blk_310_67_buf_req_0 : boolean;
  signal n_blk_310_67_buf_ack_0 : boolean;
  signal n_blk_310_67_buf_req_1 : boolean;
  signal n_blk_310_67_buf_ack_1 : boolean;
  signal phi_stmt_68_req_1 : boolean;
  signal phi_stmt_68_req_0 : boolean;
  signal phi_stmt_68_ack_0 : boolean;
  signal WPIPE_input_pipe1_169_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_169_inst_ack_1 : boolean;
  signal W_c3_166_delayed_14_0_172_inst_req_0 : boolean;
  signal W_c3_166_delayed_14_0_172_inst_ack_0 : boolean;
  signal W_c3_166_delayed_14_0_172_inst_req_1 : boolean;
  signal W_c3_166_delayed_14_0_172_inst_ack_1 : boolean;
  signal n_winr_211_72_buf_req_1 : boolean;
  signal n_winr_211_72_buf_ack_1 : boolean;
  signal phi_stmt_73_req_1 : boolean;
  signal phi_stmt_73_req_0 : boolean;
  signal phi_stmt_73_ack_0 : boolean;
  signal n_col_224_77_buf_req_0 : boolean;
  signal n_col_224_77_buf_ack_0 : boolean;
  signal n_col_224_77_buf_req_1 : boolean;
  signal n_col_224_77_buf_ack_1 : boolean;
  signal phi_stmt_78_req_0 : boolean;
  signal phi_stmt_78_req_1 : boolean;
  signal phi_stmt_78_ack_0 : boolean;
  signal n_row_236_80_buf_req_0 : boolean;
  signal n_row_236_80_buf_ack_0 : boolean;
  signal n_row_236_80_buf_req_1 : boolean;
  signal n_row_236_80_buf_ack_1 : boolean;
  signal array_obj_ref_135_index_offset_req_0 : boolean;
  signal array_obj_ref_135_index_offset_ack_0 : boolean;
  signal array_obj_ref_135_index_offset_req_1 : boolean;
  signal array_obj_ref_135_index_offset_ack_1 : boolean;
  signal addr_of_136_final_reg_req_0 : boolean;
  signal addr_of_136_final_reg_ack_0 : boolean;
  signal addr_of_136_final_reg_req_1 : boolean;
  signal addr_of_136_final_reg_ack_1 : boolean;
  signal ptr_deref_140_load_0_req_0 : boolean;
  signal ptr_deref_140_load_0_ack_0 : boolean;
  signal ptr_deref_140_load_0_req_1 : boolean;
  signal ptr_deref_140_load_0_ack_1 : boolean;
  signal slice_144_inst_req_0 : boolean;
  signal slice_144_inst_ack_0 : boolean;
  signal slice_144_inst_req_1 : boolean;
  signal slice_144_inst_ack_1 : boolean;
  signal slice_148_inst_req_0 : boolean;
  signal slice_148_inst_ack_0 : boolean;
  signal slice_148_inst_req_1 : boolean;
  signal slice_148_inst_ack_1 : boolean;
  signal slice_152_inst_req_0 : boolean;
  signal slice_152_inst_ack_0 : boolean;
  signal slice_152_inst_req_1 : boolean;
  signal slice_152_inst_ack_1 : boolean;
  signal slice_156_inst_req_0 : boolean;
  signal slice_156_inst_ack_0 : boolean;
  signal slice_156_inst_req_1 : boolean;
  signal slice_156_inst_ack_1 : boolean;
  signal W_c1_158_delayed_14_0_158_inst_req_0 : boolean;
  signal W_c1_158_delayed_14_0_158_inst_ack_0 : boolean;
  signal W_c1_158_delayed_14_0_158_inst_req_1 : boolean;
  signal W_c1_158_delayed_14_0_158_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_162_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_162_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_162_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_162_inst_ack_1 : boolean;
  signal W_c2_162_delayed_14_0_165_inst_req_0 : boolean;
  signal W_c2_162_delayed_14_0_165_inst_ack_0 : boolean;
  signal W_c2_162_delayed_14_0_165_inst_req_1 : boolean;
  signal W_c2_162_delayed_14_0_165_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_169_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_169_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_176_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_176_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_176_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_176_inst_ack_1 : boolean;
  signal W_c4_170_delayed_14_0_179_inst_req_0 : boolean;
  signal W_c4_170_delayed_14_0_179_inst_ack_0 : boolean;
  signal W_c4_170_delayed_14_0_179_inst_req_1 : boolean;
  signal W_c4_170_delayed_14_0_179_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_183_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_183_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_183_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_183_inst_ack_1 : boolean;
  signal do_while_stmt_46_branch_ack_0 : boolean;
  signal do_while_stmt_46_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 96) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= num_cont;
  num_cont_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= row1;
  row1_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= col1;
  col1_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(63 downto 48) <= rk1;
  rk1_buffer <= in_buffer_data_out(63 downto 48);
  in_buffer_data_in(79 downto 64) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(95 downto 80) <= ct;
  ct_buffer <= in_buffer_data_out(95 downto 80);
  in_buffer_data_in(tag_length + 95 downto 96) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 95 downto 96);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(207 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_34_to_assign_stmt_45/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_34_to_assign_stmt_45/$exit
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_28/$entry
      -- CP-element group 0: 	 branch_block_stmt_28/branch_block_stmt_28__entry__
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_34_to_assign_stmt_45__entry__
      -- CP-element group 0: 	 branch_block_stmt_28/assign_stmt_34_to_assign_stmt_45__exit__
      -- CP-element group 0: 	 branch_block_stmt_28/do_while_stmt_46__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	207 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_28/$exit
      -- CP-element group 1: 	 branch_block_stmt_28/branch_block_stmt_28__exit__
      -- CP-element group 1: 	 branch_block_stmt_28/do_while_stmt_46__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(207);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_28/do_while_stmt_46/$entry
      -- CP-element group 2: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46__entry__
      -- 
    access_T_CP_0_elements(2) <= access_T_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	207 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46__exit__
      -- 
    -- Element group access_T_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_28/do_while_stmt_46/loop_back
      -- 
    -- Element group access_T_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	205 
    -- CP-element group 5: 	206 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_28/do_while_stmt_46/condition_done
      -- CP-element group 5: 	 branch_block_stmt_28/do_while_stmt_46/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_28/do_while_stmt_46/loop_taken/$entry
      -- 
    access_T_CP_0_elements(5) <= access_T_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	204 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_28/do_while_stmt_46/loop_body_done
      -- 
    access_T_CP_0_elements(6) <= access_T_CP_0_elements(204);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	78 
    -- CP-element group 7: 	97 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	116 
    -- CP-element group 7: 	135 
    -- CP-element group 7: 	59 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(7) <= access_T_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	80 
    -- CP-element group 8: 	99 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	118 
    -- CP-element group 8: 	137 
    -- CP-element group 8: 	61 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(8) <= access_T_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	203 
    -- CP-element group 9: 	72 
    -- CP-element group 9: 	73 
    -- CP-element group 9: 	93 
    -- CP-element group 9: 	94 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	110 
    -- CP-element group 9: 	111 
    -- CP-element group 9: 	149 
    -- CP-element group 9: 	150 
    -- CP-element group 9: 	129 
    -- CP-element group 9: 	130 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	54 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	203 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/condition_evaluated
      -- 
    condition_evaluated_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(10), ack => do_while_stmt_46_branch_req_0); -- 
    access_T_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(203) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	93 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	110 
    -- CP-element group 11: 	129 
    -- CP-element group 11: 	53 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	74 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	112 
    -- CP-element group 11: 	131 
    -- CP-element group 11: 	55 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_sample_start__ps
      -- 
    access_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= access_T_CP_0_elements(72) & access_T_CP_0_elements(93) & access_T_CP_0_elements(15) & access_T_CP_0_elements(34) & access_T_CP_0_elements(110) & access_T_CP_0_elements(129) & access_T_CP_0_elements(53) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	95 
    -- CP-element group 12: 	75 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	113 
    -- CP-element group 12: 	132 
    -- CP-element group 12: 	56 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	204 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	72 
    -- CP-element group 12: 	93 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	110 
    -- CP-element group 12: 	129 
    -- CP-element group 12: 	53 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_sample_completed_
      -- 
    access_T_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(95) & access_T_CP_0_elements(75) & access_T_CP_0_elements(18) & access_T_CP_0_elements(37) & access_T_CP_0_elements(113) & access_T_CP_0_elements(132) & access_T_CP_0_elements(56);
      gj_access_T_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	73 
    -- CP-element group 13: 	94 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	111 
    -- CP-element group 13: 	130 
    -- CP-element group 13: 	54 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	76 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	114 
    -- CP-element group 13: 	133 
    -- CP-element group 13: 	57 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_update_start__ps
      -- 
    access_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(73) & access_T_CP_0_elements(94) & access_T_CP_0_elements(16) & access_T_CP_0_elements(35) & access_T_CP_0_elements(111) & access_T_CP_0_elements(130) & access_T_CP_0_elements(54);
      gj_access_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	77 
    -- CP-element group 14: 	96 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	115 
    -- CP-element group 14: 	134 
    -- CP-element group 14: 	58 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(77) & access_T_CP_0_elements(96) & access_T_CP_0_elements(20) & access_T_CP_0_elements(39) & access_T_CP_0_elements(115) & access_T_CP_0_elements(134) & access_T_CP_0_elements(58);
      gj_access_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_sample_start_
      -- 
    access_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	151 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_update_start_
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_sample_start__ps
      -- 
    access_T_CP_0_elements(17) <= access_T_CP_0_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_update_start__ps
      -- 
    access_T_CP_0_elements(19) <= access_T_CP_0_elements(13);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: 	151 
    -- CP-element group 20:  members (15) 
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_resized_1
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_scaled_1
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_computed_1
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_resize_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_resize_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_resize_1/index_resize_req
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_resize_1/index_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_scale_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_scale_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_scale_1/scale_rename_req
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_index_scale_1/scale_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_final_index_sum_regn_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_final_index_sum_regn_Sample/req
      -- 
    req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(20), ack => array_obj_ref_135_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_loopback_trigger
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_loopback_sample_req_ps
      -- 
    phi_stmt_48_loopback_sample_req_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_48_loopback_sample_req_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(22), ack => phi_stmt_48_req_0); -- 
    -- Element group access_T_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_entry_trigger
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_entry_sample_req_ps
      -- 
    phi_stmt_48_entry_sample_req_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_48_entry_sample_req_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(24), ack => phi_stmt_48_req_1); -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_48_phi_mux_ack_ps
      -- 
    phi_stmt_48_phi_mux_ack_50_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_48_ack_0, ack => access_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_Sample/req
      -- 
    req_63_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_63_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(26), ack => n_address_282_50_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_update_start_
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_Update/req
      -- 
    req_68_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_68_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(27), ack => n_address_282_50_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_Sample/ack
      -- 
    ack_64_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_282_50_buf_ack_0, ack => access_T_CP_0_elements(28)); -- 
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_address_50_Update/ack
      -- 
    ack_69_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_282_50_buf_ack_1, ack => access_T_CP_0_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_52_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_52_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_52_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_52_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_52_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_52_update_start_
      -- 
    -- Element group access_T_CP_0_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_52_update_completed__ps
      -- 
    access_T_CP_0_elements(32) <= access_T_CP_0_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_52_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(31), ack => access_T_CP_0_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_sample_start_
      -- 
    access_T_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	177 
    -- CP-element group 35: 	184 
    -- CP-element group 35: 	191 
    -- CP-element group 35: 	198 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_update_start_
      -- 
    access_T_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(177) & access_T_CP_0_elements(184) & access_T_CP_0_elements(191) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_sample_start__ps
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_update_start__ps
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	175 
    -- CP-element group 39: 	182 
    -- CP-element group 39: 	189 
    -- CP-element group 39: 	196 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_loopback_trigger
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_loopback_sample_req_ps
      -- 
    phi_stmt_53_loopback_sample_req_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_53_loopback_sample_req_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => phi_stmt_53_req_1); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_entry_trigger
      -- 
    access_T_CP_0_elements(42) <= access_T_CP_0_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_entry_sample_req_ps
      -- 
    phi_stmt_53_entry_sample_req_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_53_entry_sample_req_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => phi_stmt_53_req_0); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_53_phi_mux_ack_ps
      -- 
    phi_stmt_53_phi_mux_ack_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_53_ack_0, ack => access_T_CP_0_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_57_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_57_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_57_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_57_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_57_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_57_update_start_
      -- 
    -- Element group access_T_CP_0_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_57_update_completed__ps
      -- 
    access_T_CP_0_elements(47) <= access_T_CP_0_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_57_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(46), ack => access_T_CP_0_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_Sample/req
      -- 
    req_115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(49), ack => n_word_start_271_58_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_update_start_
      -- CP-element group 50: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_Update/req
      -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(50), ack => n_word_start_271_58_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_Sample/ack
      -- 
    ack_116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_271_58_buf_ack_0, ack => access_T_CP_0_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_word_start_58_Update/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_271_58_buf_ack_1, ack => access_T_CP_0_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	12 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	11 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_sample_start_
      -- 
    access_T_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	9 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	58 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	13 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_update_start_
      -- 
    access_T_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(58);
      gj_access_T_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	11 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_sample_start__ps
      -- 
    access_T_CP_0_elements(55) <= access_T_CP_0_elements(11);
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	13 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_update_start__ps
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(13);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	54 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	7 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_loopback_trigger
      -- 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(7);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_loopback_sample_req
      -- CP-element group 60: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_loopback_sample_req_ps
      -- 
    phi_stmt_59_loopback_sample_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_59_loopback_sample_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(60), ack => phi_stmt_59_req_0); -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	8 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_entry_trigger
      -- 
    access_T_CP_0_elements(61) <= access_T_CP_0_elements(8);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_entry_sample_req
      -- CP-element group 62: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_entry_sample_req_ps
      -- 
    phi_stmt_59_entry_sample_req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_59_entry_sample_req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => phi_stmt_59_req_1); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_phi_mux_ack
      -- CP-element group 63: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_59_phi_mux_ack_ps
      -- 
    phi_stmt_59_phi_mux_ack_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_59_ack_0, ack => access_T_CP_0_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_sample_start__ps
      -- CP-element group 64: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_Sample/req
      -- 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(64), ack => n_left_290_61_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_update_start__ps
      -- CP-element group 65: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_update_start_
      -- CP-element group 65: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_Update/req
      -- 
    req_156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(65), ack => n_left_290_61_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_Sample/ack
      -- 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_290_61_buf_ack_0, ack => access_T_CP_0_elements(66)); -- 
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_update_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_left_61_Update/ack
      -- 
    ack_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_290_61_buf_ack_1, ack => access_T_CP_0_elements(67)); -- 
    -- CP-element group 68:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_sample_start__ps
      -- CP-element group 68: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_Sample/req
      -- 
    req_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(68), ack => nl_start_37_62_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_update_start__ps
      -- CP-element group 69: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_update_start_
      -- CP-element group 69: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_Update/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(69), ack => nl_start_37_62_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_Sample/ack
      -- 
    ack_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_37_62_buf_ack_0, ack => access_T_CP_0_elements(70)); -- 
    -- CP-element group 71:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_update_completed__ps
      -- CP-element group 71: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_nl_start_62_Update/ack
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_37_62_buf_ack_1, ack => access_T_CP_0_elements(71)); -- 
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	9 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	12 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	11 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_sample_start_
      -- 
    access_T_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	9 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	184 
    -- CP-element group 73: 	191 
    -- CP-element group 73: 	198 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	13 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_update_start_
      -- 
    access_T_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(184) & access_T_CP_0_elements(191) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	11 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_sample_start__ps
      -- 
    access_T_CP_0_elements(74) <= access_T_CP_0_elements(11);
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	12 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	13 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_update_start__ps
      -- 
    access_T_CP_0_elements(76) <= access_T_CP_0_elements(13);
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	182 
    -- CP-element group 77: 	189 
    -- CP-element group 77: 	196 
    -- CP-element group 77: 	14 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	7 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_loopback_trigger
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(7);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_loopback_sample_req
      -- CP-element group 79: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_loopback_sample_req_ps
      -- 
    phi_stmt_63_loopback_sample_req_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_63_loopback_sample_req_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(79), ack => phi_stmt_63_req_1); -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	8 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_entry_trigger
      -- 
    access_T_CP_0_elements(80) <= access_T_CP_0_elements(8);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_entry_sample_req
      -- CP-element group 81: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_entry_sample_req_ps
      -- 
    phi_stmt_63_entry_sample_req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_63_entry_sample_req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(81), ack => phi_stmt_63_req_0); -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_phi_mux_ack
      -- CP-element group 82: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_63_phi_mux_ack_ps
      -- 
    phi_stmt_63_phi_mux_ack_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_63_ack_0, ack => access_T_CP_0_elements(82)); -- 
    -- CP-element group 83:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(84) is bound as output of CP function.
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_Sample/rr
      -- 
    rr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(85), ack => type_cast_66_inst_req_0); -- 
    access_T_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(83) & access_T_CP_0_elements(87);
      gj_access_T_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_update_start_
      -- CP-element group 86: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_Update/cr
      -- 
    cr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(86), ack => type_cast_66_inst_req_1); -- 
    access_T_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(84) & access_T_CP_0_elements(88);
      gj_access_T_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_Sample/ra
      -- 
    ra_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_66_inst_ack_0, ack => access_T_CP_0_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_update_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_66_Update/ca
      -- 
    ca_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_66_inst_ack_1, ack => access_T_CP_0_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_sample_start__ps
      -- CP-element group 89: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_Sample/req
      -- 
    req_223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(89), ack => n_blk_310_67_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_update_start__ps
      -- CP-element group 90: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_update_start_
      -- CP-element group 90: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_Update/req
      -- 
    req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(90), ack => n_blk_310_67_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_sample_completed__ps
      -- CP-element group 91: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_Sample/ack
      -- 
    ack_224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_310_67_buf_ack_0, ack => access_T_CP_0_elements(91)); -- 
    -- CP-element group 92:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_update_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_blk_67_Update/ack
      -- 
    ack_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_310_67_buf_ack_1, ack => access_T_CP_0_elements(92)); -- 
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	9 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	12 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	11 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_sample_start_
      -- 
    access_T_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	9 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	13 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_update_start_
      -- 
    access_T_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(96);
      gj_access_T_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	12 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(95) is bound as output of CP function.
    -- CP-element group 96:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	14 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	94 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	7 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_loopback_trigger
      -- 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(7);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_loopback_sample_req
      -- CP-element group 98: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_loopback_sample_req_ps
      -- 
    phi_stmt_68_loopback_sample_req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_68_loopback_sample_req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(98), ack => phi_stmt_68_req_1); -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	8 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_entry_trigger
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(8);
    -- CP-element group 100:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_entry_sample_req
      -- CP-element group 100: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_entry_sample_req_ps
      -- 
    phi_stmt_68_entry_sample_req_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_68_entry_sample_req_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(100), ack => phi_stmt_68_req_0); -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_phi_mux_ack
      -- CP-element group 101: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_68_phi_mux_ack_ps
      -- 
    phi_stmt_68_phi_mux_ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_68_ack_0, ack => access_T_CP_0_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_71_sample_start__ps
      -- CP-element group 102: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_71_sample_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_71_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_71_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_71_update_start__ps
      -- CP-element group 103: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_71_update_start_
      -- 
    -- Element group access_T_CP_0_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_71_update_completed__ps
      -- 
    access_T_CP_0_elements(104) <= access_T_CP_0_elements(105);
    -- CP-element group 105:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	104 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_71_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(103), ack => access_T_CP_0_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_sample_start__ps
      -- CP-element group 106: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_Sample/req
      -- 
    req_267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(106), ack => n_winr_211_72_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_update_start__ps
      -- CP-element group 107: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_update_start_
      -- CP-element group 107: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_Update/req
      -- 
    req_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(107), ack => n_winr_211_72_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_Sample/ack
      -- 
    ack_268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_211_72_buf_ack_0, ack => access_T_CP_0_elements(108)); -- 
    -- CP-element group 109:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_update_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_winr_72_Update/ack
      -- 
    ack_273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_211_72_buf_ack_1, ack => access_T_CP_0_elements(109)); -- 
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	9 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	12 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	11 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_sample_start_
      -- 
    access_T_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	9 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	115 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	13 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_update_start_
      -- 
    access_T_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(115);
      gj_access_T_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	11 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_sample_start__ps
      -- 
    access_T_CP_0_elements(112) <= access_T_CP_0_elements(11);
    -- CP-element group 113:  join  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	12 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(113) is bound as output of CP function.
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	13 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_update_start__ps
      -- 
    access_T_CP_0_elements(114) <= access_T_CP_0_elements(13);
    -- CP-element group 115:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	14 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	111 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	7 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_loopback_trigger
      -- 
    access_T_CP_0_elements(116) <= access_T_CP_0_elements(7);
    -- CP-element group 117:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_loopback_sample_req
      -- CP-element group 117: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_loopback_sample_req_ps
      -- 
    phi_stmt_73_loopback_sample_req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_73_loopback_sample_req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(117), ack => phi_stmt_73_req_1); -- 
    -- Element group access_T_CP_0_elements(117) is bound as output of CP function.
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	8 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_entry_trigger
      -- 
    access_T_CP_0_elements(118) <= access_T_CP_0_elements(8);
    -- CP-element group 119:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_entry_sample_req
      -- CP-element group 119: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_entry_sample_req_ps
      -- 
    phi_stmt_73_entry_sample_req_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_73_entry_sample_req_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(119), ack => phi_stmt_73_req_0); -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_phi_mux_ack
      -- CP-element group 120: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_73_phi_mux_ack_ps
      -- 
    phi_stmt_73_phi_mux_ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_73_ack_0, ack => access_T_CP_0_elements(120)); -- 
    -- CP-element group 121:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_76_sample_start__ps
      -- CP-element group 121: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_76_sample_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_76_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_76_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_76_update_start__ps
      -- CP-element group 122: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_76_update_start_
      -- 
    -- Element group access_T_CP_0_elements(122) is bound as output of CP function.
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_76_update_completed__ps
      -- 
    access_T_CP_0_elements(123) <= access_T_CP_0_elements(124);
    -- CP-element group 124:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	123 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_76_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(124) is a control-delay.
    cp_element_124_delay: control_delay_element  generic map(name => " 124_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(122), ack => access_T_CP_0_elements(124), clk => clk, reset =>reset);
    -- CP-element group 125:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_sample_start__ps
      -- CP-element group 125: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_Sample/req
      -- 
    req_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(125), ack => n_col_224_77_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_update_start__ps
      -- CP-element group 126: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_update_start_
      -- CP-element group 126: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_Update/req
      -- 
    req_316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(126), ack => n_col_224_77_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_Sample/ack
      -- 
    ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_224_77_buf_ack_0, ack => access_T_CP_0_elements(127)); -- 
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (4) 
      -- CP-element group 128: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_update_completed__ps
      -- CP-element group 128: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_col_77_Update/ack
      -- 
    ack_317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_224_77_buf_ack_1, ack => access_T_CP_0_elements(128)); -- 
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	9 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	12 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	11 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_sample_start_
      -- 
    access_T_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	9 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	134 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	13 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_update_start_
      -- 
    access_T_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	11 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_sample_start__ps
      -- 
    access_T_CP_0_elements(131) <= access_T_CP_0_elements(11);
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	12 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(132) is bound as output of CP function.
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	13 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_update_start__ps
      -- 
    access_T_CP_0_elements(133) <= access_T_CP_0_elements(13);
    -- CP-element group 134:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	14 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	130 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	7 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_loopback_trigger
      -- 
    access_T_CP_0_elements(135) <= access_T_CP_0_elements(7);
    -- CP-element group 136:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_loopback_sample_req
      -- CP-element group 136: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_loopback_sample_req_ps
      -- 
    phi_stmt_78_loopback_sample_req_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_78_loopback_sample_req_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => phi_stmt_78_req_0); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	8 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_entry_trigger
      -- 
    access_T_CP_0_elements(137) <= access_T_CP_0_elements(8);
    -- CP-element group 138:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_entry_sample_req
      -- CP-element group 138: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_entry_sample_req_ps
      -- 
    phi_stmt_78_entry_sample_req_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_78_entry_sample_req_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(138), ack => phi_stmt_78_req_1); -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_phi_mux_ack
      -- CP-element group 139: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/phi_stmt_78_phi_mux_ack_ps
      -- 
    phi_stmt_78_phi_mux_ack_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_78_ack_0, ack => access_T_CP_0_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_sample_start__ps
      -- CP-element group 140: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_Sample/req
      -- 
    req_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(140), ack => n_row_236_80_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (4) 
      -- CP-element group 141: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_update_start__ps
      -- CP-element group 141: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_update_start_
      -- CP-element group 141: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_Update/req
      -- 
    req_352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(141), ack => n_row_236_80_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_sample_completed__ps
      -- CP-element group 142: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_Sample/ack
      -- 
    ack_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_236_80_buf_ack_0, ack => access_T_CP_0_elements(142)); -- 
    -- CP-element group 143:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_update_completed__ps
      -- CP-element group 143: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/R_n_row_80_Update/ack
      -- 
    ack_353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_236_80_buf_ack_1, ack => access_T_CP_0_elements(143)); -- 
    -- CP-element group 144:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_82_sample_start__ps
      -- CP-element group 144: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_82_sample_completed__ps
      -- CP-element group 144: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_82_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_82_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_82_update_start__ps
      -- CP-element group 145: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_82_update_start_
      -- 
    -- Element group access_T_CP_0_elements(145) is bound as output of CP function.
    -- CP-element group 146:  join  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_82_update_completed__ps
      -- 
    access_T_CP_0_elements(146) <= access_T_CP_0_elements(147);
    -- CP-element group 147:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	146 
    -- CP-element group 147:  members (1) 
      -- CP-element group 147: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/type_cast_82_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(147) is a control-delay.
    cp_element_147_delay: control_delay_element  generic map(name => " 147_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(145), ack => access_T_CP_0_elements(147), clk => clk, reset =>reset);
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	152 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	153 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_request/$entry
      -- CP-element group 148: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_request/req
      -- 
    req_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(148), ack => addr_of_136_final_reg_req_0); -- 
    access_T_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(152) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	9 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	157 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	154 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_update_start_
      -- CP-element group 149: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_complete/req
      -- 
    req_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(149), ack => addr_of_136_final_reg_req_1); -- 
    access_T_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_final_index_sum_regn_update_start
      -- CP-element group 150: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_final_index_sum_regn_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_final_index_sum_regn_Update/req
      -- 
    req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => array_obj_ref_135_index_offset_req_1); -- 
    access_T_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	20 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	204 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	16 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_final_index_sum_regn_sample_complete
      -- CP-element group 151: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_final_index_sum_regn_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_final_index_sum_regn_Sample/ack
      -- 
    ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_135_index_offset_ack_0, ack => access_T_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	148 
    -- CP-element group 152:  members (8) 
      -- CP-element group 152: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_root_address_calculated
      -- CP-element group 152: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_offset_calculated
      -- CP-element group 152: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_final_index_sum_regn_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_final_index_sum_regn_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_base_plus_offset/$entry
      -- CP-element group 152: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_base_plus_offset/$exit
      -- CP-element group 152: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_base_plus_offset/sum_rename_req
      -- CP-element group 152: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/array_obj_ref_135_base_plus_offset/sum_rename_ack
      -- 
    ack_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_135_index_offset_ack_1, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_request/$exit
      -- CP-element group 153: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_request/ack
      -- 
    ack_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_136_final_reg_ack_0, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	149 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (19) 
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_complete/$exit
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/addr_of_136_complete/ack
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_word_addrgen/root_register_ack
      -- 
    ack_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_136_final_reg_ack_1, ack => access_T_CP_0_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (5) 
      -- CP-element group 155: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Sample/word_access_start/$entry
      -- CP-element group 155: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Sample/word_access_start/word_0/$entry
      -- CP-element group 155: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Sample/word_access_start/word_0/rr
      -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(155), ack => ptr_deref_140_load_0_req_0); -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(154) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	169 
    -- CP-element group 156: 	173 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	165 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_update_start_
      -- CP-element group 156: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/word_access_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/word_access_complete/word_0/$entry
      -- CP-element group 156: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/word_access_complete/word_0/cr
      -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(156), ack => ptr_deref_140_load_0_req_1); -- 
    access_T_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(169) & access_T_CP_0_elements(173) & access_T_CP_0_elements(161) & access_T_CP_0_elements(165);
      gj_access_T_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	149 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Sample/word_access_start/$exit
      -- CP-element group 157: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Sample/word_access_start/word_0/$exit
      -- CP-element group 157: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Sample/word_access_start/word_0/ra
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_140_load_0_ack_0, ack => access_T_CP_0_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	171 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	163 
    -- CP-element group 158: 	167 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/word_access_complete/$exit
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/word_access_complete/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/word_access_complete/word_0/ca
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/ptr_deref_140_Merge/$entry
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/ptr_deref_140_Merge/$exit
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/ptr_deref_140_Merge/merge_req
      -- CP-element group 158: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/ptr_deref_140_Update/ptr_deref_140_Merge/merge_ack
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_140_load_0_ack_1, ack => access_T_CP_0_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_Sample/rr
      -- 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(159), ack => slice_144_inst_req_0); -- 
    access_T_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(161);
      gj_access_T_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	180 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_update_start_
      -- CP-element group 160: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_Update/cr
      -- 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(160), ack => slice_144_inst_req_1); -- 
    access_T_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: 	156 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_Sample/ra
      -- 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_144_inst_ack_0, ack => access_T_CP_0_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	179 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_144_Update/ca
      -- 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_144_inst_ack_1, ack => access_T_CP_0_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	158 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_Sample/rr
      -- 
    rr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => slice_148_inst_req_0); -- 
    access_T_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(165);
      gj_access_T_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	187 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_update_start_
      -- CP-element group 164: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_Update/cr
      -- 
    cr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(164), ack => slice_148_inst_req_1); -- 
    access_T_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	156 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_Sample/ra
      -- 
    ra_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_148_inst_ack_0, ack => access_T_CP_0_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	186 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_148_Update/ca
      -- 
    ca_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_148_inst_ack_1, ack => access_T_CP_0_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	158 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_Sample/rr
      -- 
    rr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(167), ack => slice_152_inst_req_0); -- 
    access_T_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	194 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_update_start_
      -- CP-element group 168: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_Update/cr
      -- 
    cr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(168), ack => slice_152_inst_req_1); -- 
    access_T_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: 	156 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_Sample/ra
      -- 
    ra_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_152_inst_ack_0, ack => access_T_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	193 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_152_Update/ca
      -- 
    ca_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_152_inst_ack_1, ack => access_T_CP_0_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	158 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_Sample/rr
      -- 
    rr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(171), ack => slice_156_inst_req_0); -- 
    access_T_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(173);
      gj_access_T_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	201 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_update_start_
      -- CP-element group 172: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_Update/cr
      -- 
    cr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(172), ack => slice_156_inst_req_1); -- 
    access_T_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: 	156 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_Sample/ra
      -- 
    ra_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_156_inst_ack_0, ack => access_T_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	200 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/slice_156_Update/ca
      -- 
    ca_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_156_inst_ack_1, ack => access_T_CP_0_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	39 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_Sample/req
      -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(175), ack => W_c1_158_delayed_14_0_158_inst_req_0); -- 
    access_T_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(39) & access_T_CP_0_elements(177);
      gj_access_T_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	180 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_update_start_
      -- CP-element group 176: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_Update/req
      -- 
    req_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(176), ack => W_c1_158_delayed_14_0_158_inst_req_1); -- 
    access_T_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: 	35 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_Sample/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_158_delayed_14_0_158_inst_ack_0, ack => access_T_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_160_Update/ack
      -- 
    ack_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_158_delayed_14_0_158_inst_ack_1, ack => access_T_CP_0_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: 	162 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	202 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_Sample/req
      -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(179), ack => WPIPE_input_pipe1_162_inst_req_0); -- 
    access_T_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(178) & access_T_CP_0_elements(162) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	176 
    -- CP-element group 180: 	160 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_update_start_
      -- CP-element group 180: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_Update/req
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_162_inst_ack_0, ack => access_T_CP_0_elements(180)); -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => WPIPE_input_pipe1_162_inst_req_1); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	186 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_162_Update/ack
      -- 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_162_inst_ack_1, ack => access_T_CP_0_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	77 
    -- CP-element group 182: 	39 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_Sample/req
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => W_c2_162_delayed_14_0_165_inst_req_0); -- 
    access_T_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(77) & access_T_CP_0_elements(39) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	187 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_update_start_
      -- CP-element group 183: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_Update/req
      -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(183), ack => W_c2_162_delayed_14_0_165_inst_req_1); -- 
    access_T_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	73 
    -- CP-element group 184: 	35 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_Sample/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_162_delayed_14_0_165_inst_ack_0, ack => access_T_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_167_Update/ack
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_162_delayed_14_0_165_inst_ack_1, ack => access_T_CP_0_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	181 
    -- CP-element group 186: 	185 
    -- CP-element group 186: 	166 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_Sample/req
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(186), ack => WPIPE_input_pipe1_169_inst_req_0); -- 
    access_T_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(181) & access_T_CP_0_elements(185) & access_T_CP_0_elements(166) & access_T_CP_0_elements(188);
      gj_access_T_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	183 
    -- CP-element group 187: 	164 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_Update/req
      -- CP-element group 187: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_update_start_
      -- CP-element group 187: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_Sample/ack
      -- CP-element group 187: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_Update/$entry
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_169_inst_ack_0, ack => access_T_CP_0_elements(187)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(187), ack => WPIPE_input_pipe1_169_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	193 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_Update/ack
      -- CP-element group 188: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_169_Update/$exit
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_169_inst_ack_1, ack => access_T_CP_0_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	77 
    -- CP-element group 189: 	39 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_Sample/req
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(189), ack => W_c3_166_delayed_14_0_172_inst_req_0); -- 
    access_T_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(77) & access_T_CP_0_elements(39) & access_T_CP_0_elements(191);
      gj_access_T_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_update_start_
      -- CP-element group 190: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_Update/req
      -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(190), ack => W_c3_166_delayed_14_0_172_inst_req_1); -- 
    access_T_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: 	73 
    -- CP-element group 191: 	35 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_Sample/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_166_delayed_14_0_172_inst_ack_0, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_174_Update/ack
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_166_delayed_14_0_172_inst_ack_1, ack => access_T_CP_0_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	170 
    -- CP-element group 193: 	188 
    -- CP-element group 193: 	192 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_Sample/req
      -- 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => WPIPE_input_pipe1_176_inst_req_0); -- 
    access_T_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(170) & access_T_CP_0_elements(188) & access_T_CP_0_elements(192) & access_T_CP_0_elements(195);
      gj_access_T_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	190 
    -- CP-element group 194: 	168 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_update_start_
      -- CP-element group 194: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_Update/req
      -- 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_176_inst_ack_0, ack => access_T_CP_0_elements(194)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(194), ack => WPIPE_input_pipe1_176_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	200 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_176_Update/ack
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_176_inst_ack_1, ack => access_T_CP_0_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	77 
    -- CP-element group 196: 	39 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_Sample/req
      -- 
    req_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(196), ack => W_c4_170_delayed_14_0_179_inst_req_0); -- 
    access_T_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(77) & access_T_CP_0_elements(39) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_update_start_
      -- CP-element group 197: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_Update/req
      -- 
    req_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(197), ack => W_c4_170_delayed_14_0_179_inst_req_1); -- 
    access_T_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: 	73 
    -- CP-element group 198: 	35 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_Sample/ack
      -- 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_170_delayed_14_0_179_inst_ack_0, ack => access_T_CP_0_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/assign_stmt_181_Update/ack
      -- 
    ack_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_170_delayed_14_0_179_inst_ack_1, ack => access_T_CP_0_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	174 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	199 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_Sample/req
      -- 
    req_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(200), ack => WPIPE_input_pipe1_183_inst_req_0); -- 
    access_T_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(174) & access_T_CP_0_elements(195) & access_T_CP_0_elements(199) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	172 
    -- CP-element group 201: 	197 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_update_start_
      -- CP-element group 201: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_Update/req
      -- 
    ack_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_183_inst_ack_0, ack => access_T_CP_0_elements(201)); -- 
    req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => WPIPE_input_pipe1_183_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	179 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/WPIPE_input_pipe1_183_Update/ack
      -- 
    ack_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_183_inst_ack_1, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	9 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	10 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(203) is a control-delay.
    cp_element_203_delay: control_delay_element  generic map(name => " 203_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(9), ack => access_T_CP_0_elements(203), clk => clk, reset =>reset);
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: 	12 
    -- CP-element group 204: 	151 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	6 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_28/do_while_stmt_46/do_while_stmt_46_loop_body/$exit
      -- 
    access_T_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(202) & access_T_CP_0_elements(12) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	5 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_28/do_while_stmt_46/loop_exit/$exit
      -- CP-element group 205: 	 branch_block_stmt_28/do_while_stmt_46/loop_exit/ack
      -- 
    ack_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_46_branch_ack_0, ack => access_T_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	5 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_28/do_while_stmt_46/loop_taken/$exit
      -- CP-element group 206: 	 branch_block_stmt_28/do_while_stmt_46/loop_taken/ack
      -- 
    ack_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_46_branch_ack_1, ack => access_T_CP_0_elements(206)); -- 
    -- CP-element group 207:  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	3 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	1 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_28/do_while_stmt_46/$exit
      -- 
    access_T_CP_0_elements(207) <= access_T_CP_0_elements(3);
    access_T_do_while_stmt_46_terminator_636: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_46_terminator_636", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(6),loop_continue => access_T_CP_0_elements(206),loop_terminate => access_T_CP_0_elements(205),loop_back => access_T_CP_0_elements(4),loop_exit => access_T_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_48_phi_seq_78_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(21);
      access_T_CP_0_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(28);
      access_T_CP_0_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(29);
      access_T_CP_0_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(23);
      access_T_CP_0_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(30);
      access_T_CP_0_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(32);
      access_T_CP_0_elements(24) <= phi_mux_reqs(1);
      phi_stmt_48_phi_seq_78 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_48_phi_seq_78") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(17), 
          phi_sample_ack => access_T_CP_0_elements(18), 
          phi_update_req => access_T_CP_0_elements(19), 
          phi_update_ack => access_T_CP_0_elements(20), 
          phi_mux_ack => access_T_CP_0_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_53_phi_seq_122_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(42);
      access_T_CP_0_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(45);
      access_T_CP_0_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(40);
      access_T_CP_0_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(51);
      access_T_CP_0_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(52);
      access_T_CP_0_elements(41) <= phi_mux_reqs(1);
      phi_stmt_53_phi_seq_122 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_53_phi_seq_122") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(36), 
          phi_sample_ack => access_T_CP_0_elements(37), 
          phi_update_req => access_T_CP_0_elements(38), 
          phi_update_ack => access_T_CP_0_elements(39), 
          phi_mux_ack => access_T_CP_0_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_59_phi_seq_176_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(59);
      access_T_CP_0_elements(64)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(66);
      access_T_CP_0_elements(65)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(67);
      access_T_CP_0_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(61);
      access_T_CP_0_elements(68)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(70);
      access_T_CP_0_elements(69)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(71);
      access_T_CP_0_elements(62) <= phi_mux_reqs(1);
      phi_stmt_59_phi_seq_176 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_59_phi_seq_176") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(55), 
          phi_sample_ack => access_T_CP_0_elements(56), 
          phi_update_req => access_T_CP_0_elements(57), 
          phi_update_ack => access_T_CP_0_elements(58), 
          phi_mux_ack => access_T_CP_0_elements(63), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_63_phi_seq_230_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(80);
      access_T_CP_0_elements(83)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(87);
      access_T_CP_0_elements(84)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(88);
      access_T_CP_0_elements(81) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(78);
      access_T_CP_0_elements(89)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(91);
      access_T_CP_0_elements(90)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(92);
      access_T_CP_0_elements(79) <= phi_mux_reqs(1);
      phi_stmt_63_phi_seq_230 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_63_phi_seq_230") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(74), 
          phi_sample_ack => access_T_CP_0_elements(75), 
          phi_update_req => access_T_CP_0_elements(76), 
          phi_update_ack => access_T_CP_0_elements(77), 
          phi_mux_ack => access_T_CP_0_elements(82), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_68_phi_seq_274_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(99);
      access_T_CP_0_elements(102)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(102);
      access_T_CP_0_elements(103)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(104);
      access_T_CP_0_elements(100) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(97);
      access_T_CP_0_elements(106)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(108);
      access_T_CP_0_elements(107)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(109);
      access_T_CP_0_elements(98) <= phi_mux_reqs(1);
      phi_stmt_68_phi_seq_274 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_68_phi_seq_274") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(11), 
          phi_sample_ack => access_T_CP_0_elements(95), 
          phi_update_req => access_T_CP_0_elements(13), 
          phi_update_ack => access_T_CP_0_elements(96), 
          phi_mux_ack => access_T_CP_0_elements(101), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_73_phi_seq_318_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(118);
      access_T_CP_0_elements(121)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(121);
      access_T_CP_0_elements(122)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(123);
      access_T_CP_0_elements(119) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(116);
      access_T_CP_0_elements(125)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(127);
      access_T_CP_0_elements(126)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(128);
      access_T_CP_0_elements(117) <= phi_mux_reqs(1);
      phi_stmt_73_phi_seq_318 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_73_phi_seq_318") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(112), 
          phi_sample_ack => access_T_CP_0_elements(113), 
          phi_update_req => access_T_CP_0_elements(114), 
          phi_update_ack => access_T_CP_0_elements(115), 
          phi_mux_ack => access_T_CP_0_elements(120), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_78_phi_seq_362_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(140)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(142);
      access_T_CP_0_elements(141)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(143);
      access_T_CP_0_elements(136) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(137);
      access_T_CP_0_elements(144)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(144);
      access_T_CP_0_elements(145)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(146);
      access_T_CP_0_elements(138) <= phi_mux_reqs(1);
      phi_stmt_78_phi_seq_362 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_78_phi_seq_362") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(131), 
          phi_sample_ack => access_T_CP_0_elements(132), 
          phi_update_req => access_T_CP_0_elements(133), 
          phi_update_ack => access_T_CP_0_elements(134), 
          phi_mux_ack => access_T_CP_0_elements(139), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(7);
        preds(1)  <= access_T_CP_0_elements(8);
        entry_tmerge_30 : transition_merge -- 
          generic map(name => " entry_tmerge_30")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_127_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_207_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_220_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_233_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_243_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_295_wire : std_logic_vector(15 downto 0);
    signal ADD_u64_u64_280_wire : std_logic_vector(63 downto 0);
    signal AND_u1_u1_109_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_116_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_215_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_229_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_230_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_96_wire : std_logic_vector(0 downto 0);
    signal AND_u32_u32_262_wire : std_logic_vector(31 downto 0);
    signal EQ_u2_u1_105_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_112_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_119_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_92_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_99_wire : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_276_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_242_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_244_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_32_wire : std_logic_vector(15 downto 0);
    signal MUL_u32_u32_251_wire : std_logic_vector(31 downto 0);
    signal MUX_208_wire : std_logic_vector(15 downto 0);
    signal MUX_221_wire : std_logic_vector(15 downto 0);
    signal MUX_302_wire : std_logic_vector(15 downto 0);
    signal MUX_308_wire : std_logic_vector(15 downto 0);
    signal NEQ_u16_u1_314_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_120_wire : std_logic_vector(0 downto 0);
    signal R_address_134_resized : std_logic_vector(13 downto 0);
    signal R_address_134_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_288_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_300_wire : std_logic_vector(15 downto 0);
    signal UGT_u16_u1_108_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_115_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_297_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_95_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_305_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_41_wire : std_logic_vector(0 downto 0);
    signal address_48 : std_logic_vector(63 downto 0);
    signal array_obj_ref_135_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_135_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_135_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_135_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_135_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_135_root_address : std_logic_vector(13 downto 0);
    signal c1_158_delayed_14_0_160 : std_logic_vector(0 downto 0);
    signal c1_88 : std_logic_vector(0 downto 0);
    signal c2_101 : std_logic_vector(0 downto 0);
    signal c2_162_delayed_14_0_167 : std_logic_vector(0 downto 0);
    signal c3_122 : std_logic_vector(0 downto 0);
    signal c3_166_delayed_14_0_174 : std_logic_vector(0 downto 0);
    signal c4_130 : std_logic_vector(0 downto 0);
    signal c4_170_delayed_14_0_181 : std_logic_vector(0 downto 0);
    signal col_73 : std_logic_vector(15 downto 0);
    signal col_done_200 : std_logic_vector(0 downto 0);
    signal fetch_addr_137 : std_logic_vector(31 downto 0);
    signal flag1_190 : std_logic_vector(0 downto 0);
    signal fn_blk_45 : std_logic_vector(15 downto 0);
    signal konst_104_wire_constant : std_logic_vector(1 downto 0);
    signal konst_107_wire_constant : std_logic_vector(15 downto 0);
    signal konst_111_wire_constant : std_logic_vector(1 downto 0);
    signal konst_114_wire_constant : std_logic_vector(15 downto 0);
    signal konst_118_wire_constant : std_logic_vector(1 downto 0);
    signal konst_128_wire_constant : std_logic_vector(15 downto 0);
    signal konst_204_wire_constant : std_logic_vector(15 downto 0);
    signal konst_206_wire_constant : std_logic_vector(15 downto 0);
    signal konst_217_wire_constant : std_logic_vector(15 downto 0);
    signal konst_219_wire_constant : std_logic_vector(15 downto 0);
    signal konst_232_wire_constant : std_logic_vector(15 downto 0);
    signal konst_261_wire_constant : std_logic_vector(31 downto 0);
    signal konst_269_wire_constant : std_logic_vector(1 downto 0);
    signal konst_275_wire_constant : std_logic_vector(31 downto 0);
    signal konst_279_wire_constant : std_logic_vector(63 downto 0);
    signal konst_296_wire_constant : std_logic_vector(15 downto 0);
    signal konst_298_wire_constant : std_logic_vector(15 downto 0);
    signal konst_304_wire_constant : std_logic_vector(15 downto 0);
    signal konst_307_wire_constant : std_logic_vector(15 downto 0);
    signal konst_40_wire_constant : std_logic_vector(15 downto 0);
    signal konst_43_wire_constant : std_logic_vector(15 downto 0);
    signal konst_86_wire_constant : std_logic_vector(1 downto 0);
    signal konst_91_wire_constant : std_logic_vector(1 downto 0);
    signal konst_94_wire_constant : std_logic_vector(15 downto 0);
    signal konst_98_wire_constant : std_logic_vector(1 downto 0);
    signal m_factor_34 : std_logic_vector(31 downto 0);
    signal n_address_282 : std_logic_vector(63 downto 0);
    signal n_address_282_50_buffered : std_logic_vector(63 downto 0);
    signal n_blk_310 : std_logic_vector(15 downto 0);
    signal n_blk_310_67_buffered : std_logic_vector(15 downto 0);
    signal n_col_224 : std_logic_vector(15 downto 0);
    signal n_col_224_77_buffered : std_logic_vector(15 downto 0);
    signal n_left_290 : std_logic_vector(15 downto 0);
    signal n_left_290_61_buffered : std_logic_vector(15 downto 0);
    signal n_row_236 : std_logic_vector(15 downto 0);
    signal n_row_236_80_buffered : std_logic_vector(15 downto 0);
    signal n_winr_211 : std_logic_vector(15 downto 0);
    signal n_winr_211_72_buffered : std_logic_vector(15 downto 0);
    signal n_word_start_271 : std_logic_vector(1 downto 0);
    signal n_word_start_271_58_buffered : std_logic_vector(1 downto 0);
    signal na1_246 : std_logic_vector(31 downto 0);
    signal na2_253 : std_logic_vector(31 downto 0);
    signal na3_258 : std_logic_vector(31 downto 0);
    signal na4_264 : std_logic_vector(15 downto 0);
    signal nl_start_37 : std_logic_vector(15 downto 0);
    signal nl_start_37_62_buffered : std_logic_vector(15 downto 0);
    signal num_blk_63 : std_logic_vector(15 downto 0);
    signal num_left_59 : std_logic_vector(15 downto 0);
    signal ptr_deref_140_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_140_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_140_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_140_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_140_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_78 : std_logic_vector(15 downto 0);
    signal type_cast_126_wire : std_logic_vector(15 downto 0);
    signal type_cast_250_wire : std_logic_vector(31 downto 0);
    signal type_cast_268_wire : std_logic_vector(1 downto 0);
    signal type_cast_277_wire : std_logic_vector(63 downto 0);
    signal type_cast_52_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_57_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_66_wire : std_logic_vector(15 downto 0);
    signal type_cast_71_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_76_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_82_wire_constant : std_logic_vector(15 downto 0);
    signal w1_145 : std_logic_vector(15 downto 0);
    signal w2_149 : std_logic_vector(15 downto 0);
    signal w3_153 : std_logic_vector(15 downto 0);
    signal w4_157 : std_logic_vector(15 downto 0);
    signal winr_68 : std_logic_vector(15 downto 0);
    signal winr_done_195 : std_logic_vector(0 downto 0);
    signal word_read_141 : std_logic_vector(63 downto 0);
    signal word_start_53 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_135_constant_part_of_offset <= "00000000000000";
    array_obj_ref_135_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_135_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_135_resized_base_address <= "00000000000000";
    konst_104_wire_constant <= "00";
    konst_107_wire_constant <= "0000000000000010";
    konst_111_wire_constant <= "01";
    konst_114_wire_constant <= "0000000000000001";
    konst_118_wire_constant <= "10";
    konst_128_wire_constant <= "0000000000000011";
    konst_204_wire_constant <= "0000000000000000";
    konst_206_wire_constant <= "0000000000000001";
    konst_217_wire_constant <= "0000000000000000";
    konst_219_wire_constant <= "0000000000000001";
    konst_232_wire_constant <= "0000000000000001";
    konst_261_wire_constant <= "00000000000000000000000000000011";
    konst_269_wire_constant <= "00";
    konst_275_wire_constant <= "00000000000000000000000000000010";
    konst_279_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_296_wire_constant <= "0000000000000100";
    konst_298_wire_constant <= "0000000000000100";
    konst_304_wire_constant <= "0000000000000100";
    konst_307_wire_constant <= "0000000000000100";
    konst_40_wire_constant <= "0000000000000100";
    konst_43_wire_constant <= "0000000000000100";
    konst_86_wire_constant <= "00";
    konst_91_wire_constant <= "00";
    konst_94_wire_constant <= "0000000000000001";
    konst_98_wire_constant <= "01";
    ptr_deref_140_word_offset_0 <= "00000000000000";
    type_cast_52_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_57_wire_constant <= "00";
    type_cast_71_wire_constant <= "0000000000000000";
    type_cast_76_wire_constant <= "0000000000000000";
    type_cast_82_wire_constant <= "0000000000000000";
    phi_stmt_48: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address_282_50_buffered & type_cast_52_wire_constant;
      req <= phi_stmt_48_req_0 & phi_stmt_48_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_48",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_48_ack_0,
          idata => idata,
          odata => address_48,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_48
    phi_stmt_53: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_57_wire_constant & n_word_start_271_58_buffered;
      req <= phi_stmt_53_req_0 & phi_stmt_53_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_53",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_53_ack_0,
          idata => idata,
          odata => word_start_53,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_53
    phi_stmt_59: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_left_290_61_buffered & nl_start_37_62_buffered;
      req <= phi_stmt_59_req_0 & phi_stmt_59_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_59",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_59_ack_0,
          idata => idata,
          odata => num_left_59,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_59
    phi_stmt_63: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_66_wire & n_blk_310_67_buffered;
      req <= phi_stmt_63_req_0 & phi_stmt_63_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_63",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_63_ack_0,
          idata => idata,
          odata => num_blk_63,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_63
    phi_stmt_68: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_71_wire_constant & n_winr_211_72_buffered;
      req <= phi_stmt_68_req_0 & phi_stmt_68_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_68",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_68_ack_0,
          idata => idata,
          odata => winr_68,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_68
    phi_stmt_73: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_76_wire_constant & n_col_224_77_buffered;
      req <= phi_stmt_73_req_0 & phi_stmt_73_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_73",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_73_ack_0,
          idata => idata,
          odata => col_73,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_73
    phi_stmt_78: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_row_236_80_buffered & type_cast_82_wire_constant;
      req <= phi_stmt_78_req_0 & phi_stmt_78_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_78",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_78_ack_0,
          idata => idata,
          odata => row_78,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_78
    -- flow-through select operator MUX_208_inst
    MUX_208_wire <= konst_204_wire_constant when (winr_done_195(0) /=  '0') else ADD_u16_u16_207_wire;
    -- flow-through select operator MUX_210_inst
    n_winr_211 <= MUX_208_wire when (flag1_190(0) /=  '0') else winr_68;
    -- flow-through select operator MUX_221_inst
    MUX_221_wire <= konst_217_wire_constant when (col_done_200(0) /=  '0') else ADD_u16_u16_220_wire;
    -- flow-through select operator MUX_223_inst
    n_col_224 <= MUX_221_wire when (AND_u1_u1_215_wire(0) /=  '0') else col_73;
    -- flow-through select operator MUX_235_inst
    n_row_236 <= ADD_u16_u16_233_wire when (AND_u1_u1_230_wire(0) /=  '0') else row_78;
    -- flow-through select operator MUX_270_inst
    n_word_start_271 <= type_cast_268_wire when (flag1_190(0) /=  '0') else konst_269_wire_constant;
    -- flow-through select operator MUX_281_inst
    n_address_282 <= type_cast_277_wire when (flag1_190(0) /=  '0') else ADD_u64_u64_280_wire;
    -- flow-through select operator MUX_289_inst
    n_left_290 <= nl_start_37 when (flag1_190(0) /=  '0') else SUB_u16_u16_288_wire;
    -- flow-through select operator MUX_302_inst
    MUX_302_wire <= SUB_u16_u16_300_wire when (UGT_u16_u1_297_wire(0) /=  '0') else fn_blk_45;
    -- flow-through select operator MUX_308_inst
    MUX_308_wire <= n_left_290 when (ULT_u16_u1_305_wire(0) /=  '0') else konst_307_wire_constant;
    -- flow-through select operator MUX_309_inst
    n_blk_310 <= MUX_302_wire when (flag1_190(0) /=  '0') else MUX_308_wire;
    -- flow-through select operator MUX_44_inst
    fn_blk_45 <= num_cont_buffer when (ULT_u16_u1_41_wire(0) /=  '0') else konst_43_wire_constant;
    slice_144_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_144_inst_req_0;
      slice_144_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_144_inst_req_1;
      slice_144_inst_ack_1<= update_ack(0);
      slice_144_inst: SliceSplitProtocol generic map(name => "slice_144_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_141, dout => w1_145, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_148_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_148_inst_req_0;
      slice_148_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_148_inst_req_1;
      slice_148_inst_ack_1<= update_ack(0);
      slice_148_inst: SliceSplitProtocol generic map(name => "slice_148_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_141, dout => w2_149, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_152_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_152_inst_req_0;
      slice_152_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_152_inst_req_1;
      slice_152_inst_ack_1<= update_ack(0);
      slice_152_inst: SliceSplitProtocol generic map(name => "slice_152_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_141, dout => w3_153, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_156_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_156_inst_req_0;
      slice_156_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_156_inst_req_1;
      slice_156_inst_ack_1<= update_ack(0);
      slice_156_inst: SliceSplitProtocol generic map(name => "slice_156_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_141, dout => w4_157, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_c1_158_delayed_14_0_158_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c1_158_delayed_14_0_158_inst_req_0;
      W_c1_158_delayed_14_0_158_inst_ack_0<= wack(0);
      rreq(0) <= W_c1_158_delayed_14_0_158_inst_req_1;
      W_c1_158_delayed_14_0_158_inst_ack_1<= rack(0);
      W_c1_158_delayed_14_0_158_inst : InterlockBuffer generic map ( -- 
        name => "W_c1_158_delayed_14_0_158_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c1_88,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c1_158_delayed_14_0_160,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c2_162_delayed_14_0_165_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c2_162_delayed_14_0_165_inst_req_0;
      W_c2_162_delayed_14_0_165_inst_ack_0<= wack(0);
      rreq(0) <= W_c2_162_delayed_14_0_165_inst_req_1;
      W_c2_162_delayed_14_0_165_inst_ack_1<= rack(0);
      W_c2_162_delayed_14_0_165_inst : InterlockBuffer generic map ( -- 
        name => "W_c2_162_delayed_14_0_165_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c2_101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c2_162_delayed_14_0_167,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c3_166_delayed_14_0_172_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c3_166_delayed_14_0_172_inst_req_0;
      W_c3_166_delayed_14_0_172_inst_ack_0<= wack(0);
      rreq(0) <= W_c3_166_delayed_14_0_172_inst_req_1;
      W_c3_166_delayed_14_0_172_inst_ack_1<= rack(0);
      W_c3_166_delayed_14_0_172_inst : InterlockBuffer generic map ( -- 
        name => "W_c3_166_delayed_14_0_172_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c3_122,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c3_166_delayed_14_0_174,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c4_170_delayed_14_0_179_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c4_170_delayed_14_0_179_inst_req_0;
      W_c4_170_delayed_14_0_179_inst_ack_0<= wack(0);
      rreq(0) <= W_c4_170_delayed_14_0_179_inst_req_1;
      W_c4_170_delayed_14_0_179_inst_ack_1<= rack(0);
      W_c4_170_delayed_14_0_179_inst : InterlockBuffer generic map ( -- 
        name => "W_c4_170_delayed_14_0_179_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c4_130,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c4_170_delayed_14_0_181,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_nl_start_35_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := num_cont_buffer(15 downto 0);
      nl_start_37 <= tmp_var; -- 
    end process;
    addr_of_136_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_136_final_reg_req_0;
      addr_of_136_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_136_final_reg_req_1;
      addr_of_136_final_reg_ack_1<= rack(0);
      addr_of_136_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_136_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_135_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_137,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address_282_50_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address_282_50_buf_req_0;
      n_address_282_50_buf_ack_0<= wack(0);
      rreq(0) <= n_address_282_50_buf_req_1;
      n_address_282_50_buf_ack_1<= rack(0);
      n_address_282_50_buf : InterlockBuffer generic map ( -- 
        name => "n_address_282_50_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address_282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address_282_50_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_blk_310_67_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_blk_310_67_buf_req_0;
      n_blk_310_67_buf_ack_0<= wack(0);
      rreq(0) <= n_blk_310_67_buf_req_1;
      n_blk_310_67_buf_ack_1<= rack(0);
      n_blk_310_67_buf : InterlockBuffer generic map ( -- 
        name => "n_blk_310_67_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_blk_310,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_blk_310_67_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_224_77_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_224_77_buf_req_0;
      n_col_224_77_buf_ack_0<= wack(0);
      rreq(0) <= n_col_224_77_buf_req_1;
      n_col_224_77_buf_ack_1<= rack(0);
      n_col_224_77_buf : InterlockBuffer generic map ( -- 
        name => "n_col_224_77_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_224,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_224_77_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_left_290_61_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_left_290_61_buf_req_0;
      n_left_290_61_buf_ack_0<= wack(0);
      rreq(0) <= n_left_290_61_buf_req_1;
      n_left_290_61_buf_ack_1<= rack(0);
      n_left_290_61_buf : InterlockBuffer generic map ( -- 
        name => "n_left_290_61_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_left_290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_left_290_61_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_236_80_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_236_80_buf_req_0;
      n_row_236_80_buf_ack_0<= wack(0);
      rreq(0) <= n_row_236_80_buf_req_1;
      n_row_236_80_buf_ack_1<= rack(0);
      n_row_236_80_buf : InterlockBuffer generic map ( -- 
        name => "n_row_236_80_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_236,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_236_80_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_winr_211_72_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_winr_211_72_buf_req_0;
      n_winr_211_72_buf_ack_0<= wack(0);
      rreq(0) <= n_winr_211_72_buf_req_1;
      n_winr_211_72_buf_ack_1<= rack(0);
      n_winr_211_72_buf : InterlockBuffer generic map ( -- 
        name => "n_winr_211_72_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_winr_211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_winr_211_72_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_word_start_271_58_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_word_start_271_58_buf_req_0;
      n_word_start_271_58_buf_ack_0<= wack(0);
      rreq(0) <= n_word_start_271_58_buf_req_1;
      n_word_start_271_58_buf_ack_1<= rack(0);
      n_word_start_271_58_buf : InterlockBuffer generic map ( -- 
        name => "n_word_start_271_58_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_word_start_271,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_word_start_271_58_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nl_start_37_62_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nl_start_37_62_buf_req_0;
      nl_start_37_62_buf_ack_0<= wack(0);
      rreq(0) <= nl_start_37_62_buf_req_1;
      nl_start_37_62_buf_ack_1<= rack(0);
      nl_start_37_62_buf : InterlockBuffer generic map ( -- 
        name => "nl_start_37_62_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nl_start_37,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nl_start_37_62_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_126_inst
    process(word_start_53) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := word_start_53(1 downto 0);
      type_cast_126_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_245_inst
    process(MUL_u16_u16_244_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_244_wire(15 downto 0);
      na1_246 <= tmp_var; -- 
    end process;
    -- interlock type_cast_250_inst
    process(n_winr_211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_winr_211(15 downto 0);
      type_cast_250_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_252_inst
    process(MUL_u32_u32_251_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := MUL_u32_u32_251_wire(31 downto 0);
      na2_253 <= tmp_var; -- 
    end process;
    -- interlock type_cast_263_inst
    process(AND_u32_u32_262_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := AND_u32_u32_262_wire(15 downto 0);
      na4_264 <= tmp_var; -- 
    end process;
    -- interlock type_cast_268_inst
    process(na4_264) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := na4_264(1 downto 0);
      type_cast_268_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_277_inst
    process(LSHR_u32_u32_276_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_276_wire(31 downto 0);
      type_cast_277_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_33_inst
    process(MUL_u16_u16_32_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_32_wire(15 downto 0);
      m_factor_34 <= tmp_var; -- 
    end process;
    type_cast_66_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_66_inst_req_0;
      type_cast_66_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_66_inst_req_1;
      type_cast_66_inst_ack_1<= rack(0);
      type_cast_66_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_66_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_blk_45,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_66_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_135_index_1_rename
    process(R_address_134_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_134_resized;
      ov(13 downto 0) := iv;
      R_address_134_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_135_index_1_resize
    process(address_48) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_48;
      ov := iv(13 downto 0);
      R_address_134_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_135_root_address_inst
    process(array_obj_ref_135_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_135_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_135_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_140_addr_0
    process(ptr_deref_140_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_140_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_140_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_140_base_resize
    process(fetch_addr_137) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_137;
      ov := iv(13 downto 0);
      ptr_deref_140_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_140_gather_scatter
    process(ptr_deref_140_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_140_data_0;
      ov(63 downto 0) := iv;
      word_read_141 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_140_root_address_inst
    process(ptr_deref_140_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_140_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_140_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_46_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NEQ_u16_u1_314_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_46_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_46_branch_req_0,
          ack0 => do_while_stmt_46_branch_ack_0,
          ack1 => do_while_stmt_46_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_127_inst
    process(num_blk_63, type_cast_126_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_blk_63, type_cast_126_wire, tmp_var);
      ADD_u16_u16_127_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_207_inst
    process(winr_68) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(winr_68, konst_206_wire_constant, tmp_var);
      ADD_u16_u16_207_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_220_inst
    process(col_73) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_73, konst_219_wire_constant, tmp_var);
      ADD_u16_u16_220_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_233_inst
    process(row_78) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_78, konst_232_wire_constant, tmp_var);
      ADD_u16_u16_233_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_243_inst
    process(n_col_224, MUL_u16_u16_242_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(n_col_224, MUL_u16_u16_242_wire, tmp_var);
      ADD_u16_u16_243_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_295_inst
    process(fn_blk_45, na4_264) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(fn_blk_45, na4_264, tmp_var);
      ADD_u16_u16_295_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_257_inst
    process(na1_246, na2_253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(na1_246, na2_253, tmp_var);
      na3_258 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_280_inst
    process(address_48) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_48, konst_279_wire_constant, tmp_var);
      ADD_u64_u64_280_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_109_inst
    process(EQ_u2_u1_105_wire, UGT_u16_u1_108_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_105_wire, UGT_u16_u1_108_wire, tmp_var);
      AND_u1_u1_109_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_116_inst
    process(EQ_u2_u1_112_wire, UGT_u16_u1_115_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_112_wire, UGT_u16_u1_115_wire, tmp_var);
      AND_u1_u1_116_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_215_inst
    process(winr_done_195, flag1_190) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_195, flag1_190, tmp_var);
      AND_u1_u1_215_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_229_inst
    process(col_done_200, flag1_190) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_200, flag1_190, tmp_var);
      AND_u1_u1_229_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_230_inst
    process(winr_done_195, AND_u1_u1_229_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_195, AND_u1_u1_229_wire, tmp_var);
      AND_u1_u1_230_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_96_inst
    process(EQ_u2_u1_92_wire, UGT_u16_u1_95_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_92_wire, UGT_u16_u1_95_wire, tmp_var);
      AND_u1_u1_96_wire <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_262_inst
    process(na3_258) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(na3_258, konst_261_wire_constant, tmp_var);
      AND_u32_u32_262_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_189_inst
    process(num_left_59, num_blk_63) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_left_59, num_blk_63, tmp_var);
      flag1_190 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_194_inst
    process(winr_68, rk1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(winr_68, rk1_buffer, tmp_var);
      winr_done_195 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_199_inst
    process(col_73, col1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_73, col1_buffer, tmp_var);
      col_done_200 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_105_inst
    process(word_start_53) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_53, konst_104_wire_constant, tmp_var);
      EQ_u2_u1_105_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_112_inst
    process(word_start_53) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_53, konst_111_wire_constant, tmp_var);
      EQ_u2_u1_112_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_119_inst
    process(word_start_53) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_53, konst_118_wire_constant, tmp_var);
      EQ_u2_u1_119_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_87_inst
    process(word_start_53) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_53, konst_86_wire_constant, tmp_var);
      c1_88 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_92_inst
    process(word_start_53) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_53, konst_91_wire_constant, tmp_var);
      EQ_u2_u1_92_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_99_inst
    process(word_start_53) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_53, konst_98_wire_constant, tmp_var);
      EQ_u2_u1_99_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_276_inst
    process(na3_258) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(na3_258, konst_275_wire_constant, tmp_var);
      LSHR_u32_u32_276_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_242_inst
    process(ct_buffer, n_row_236) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, n_row_236, tmp_var);
      MUL_u16_u16_242_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_244_inst
    process(chl_in_buffer, ADD_u16_u16_243_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_in_buffer, ADD_u16_u16_243_wire, tmp_var);
      MUL_u16_u16_244_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_32_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_32_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_251_inst
    process(m_factor_34, type_cast_250_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(m_factor_34, type_cast_250_wire, tmp_var);
      MUL_u32_u32_251_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u16_u1_314_inst
    process(n_row_236, row1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(n_row_236, row1_buffer, tmp_var);
      NEQ_u16_u1_314_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_100_inst
    process(AND_u1_u1_96_wire, EQ_u2_u1_99_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_96_wire, EQ_u2_u1_99_wire, tmp_var);
      c2_101 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_120_inst
    process(AND_u1_u1_116_wire, EQ_u2_u1_119_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_116_wire, EQ_u2_u1_119_wire, tmp_var);
      OR_u1_u1_120_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_121_inst
    process(AND_u1_u1_109_wire, OR_u1_u1_120_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_109_wire, OR_u1_u1_120_wire, tmp_var);
      c3_122 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_288_inst
    process(num_left_59, num_blk_63) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(num_left_59, num_blk_63, tmp_var);
      SUB_u16_u16_288_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_300_inst
    process(konst_298_wire_constant, na4_264) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_298_wire_constant, na4_264, tmp_var);
      SUB_u16_u16_300_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_108_inst
    process(num_blk_63) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_63, konst_107_wire_constant, tmp_var);
      UGT_u16_u1_108_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_115_inst
    process(num_blk_63) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_63, konst_114_wire_constant, tmp_var);
      UGT_u16_u1_115_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_129_inst
    process(ADD_u16_u16_127_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_127_wire, konst_128_wire_constant, tmp_var);
      c4_130 <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_297_inst
    process(ADD_u16_u16_295_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_295_wire, konst_296_wire_constant, tmp_var);
      UGT_u16_u1_297_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_95_inst
    process(num_blk_63) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_63, konst_94_wire_constant, tmp_var);
      UGT_u16_u1_95_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_305_inst
    process(n_left_290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_left_290, konst_304_wire_constant, tmp_var);
      ULT_u16_u1_305_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_41_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(num_cont_buffer, konst_40_wire_constant, tmp_var);
      ULT_u16_u1_41_wire <= tmp_var; --
    end process;
    -- shared split operator group (42) : array_obj_ref_135_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_134_scaled;
      array_obj_ref_135_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_135_index_offset_req_0;
      array_obj_ref_135_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_135_index_offset_req_1;
      array_obj_ref_135_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared load operator group (0) : ptr_deref_140_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_140_load_0_req_0;
      ptr_deref_140_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_140_load_0_req_1;
      ptr_deref_140_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_140_word_address_0;
      ptr_deref_140_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_169_inst WPIPE_input_pipe1_162_inst WPIPE_input_pipe1_183_inst WPIPE_input_pipe1_176_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe1_169_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe1_162_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe1_183_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe1_176_inst_req_0;
      WPIPE_input_pipe1_169_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe1_162_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe1_183_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe1_176_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe1_169_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe1_162_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe1_183_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe1_176_inst_req_1;
      WPIPE_input_pipe1_169_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe1_162_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe1_183_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe1_176_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= c3_166_delayed_14_0_174(0);
      guard_vector(1)  <= c4_170_delayed_14_0_181(0);
      guard_vector(2)  <= c1_158_delayed_14_0_160(0);
      guard_vector(3)  <= c2_162_delayed_14_0_167(0);
      data_in <= w2_149 & w1_145 & w4_157 & w3_153;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(95 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(135 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_1129_start: Boolean;
  signal convolution3D_CP_1129_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      pp : in  std_logic_vector(7 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_632_inst_req_0 : boolean;
  signal type_cast_649_inst_req_1 : boolean;
  signal type_cast_678_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_645_inst_req_1 : boolean;
  signal type_cast_561_inst_ack_0 : boolean;
  signal type_cast_524_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_532_inst_req_1 : boolean;
  signal type_cast_624_inst_ack_0 : boolean;
  signal type_cast_536_inst_ack_1 : boolean;
  signal type_cast_636_inst_req_0 : boolean;
  signal ptr_deref_1096_store_0_ack_0 : boolean;
  signal type_cast_624_inst_req_0 : boolean;
  signal type_cast_536_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_520_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_520_inst_req_0 : boolean;
  signal type_cast_574_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_532_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_ack_0 : boolean;
  signal type_cast_561_inst_req_0 : boolean;
  signal type_cast_561_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_req_1 : boolean;
  signal type_cast_561_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_620_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_req_1 : boolean;
  signal type_cast_586_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_545_inst_req_1 : boolean;
  signal type_cast_549_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_req_0 : boolean;
  signal type_cast_586_inst_req_0 : boolean;
  signal type_cast_574_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_645_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_620_inst_ack_0 : boolean;
  signal type_cast_599_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_545_inst_ack_1 : boolean;
  signal type_cast_658_inst_req_0 : boolean;
  signal type_cast_549_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_532_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_520_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_532_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_595_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_520_inst_req_1 : boolean;
  signal type_cast_599_inst_ack_0 : boolean;
  signal type_cast_649_inst_ack_1 : boolean;
  signal type_cast_611_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_ack_0 : boolean;
  signal type_cast_586_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_ack_1 : boolean;
  signal type_cast_636_inst_ack_0 : boolean;
  signal type_cast_658_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_545_inst_req_0 : boolean;
  signal type_cast_662_inst_req_1 : boolean;
  signal phi_stmt_1427_ack_0 : boolean;
  signal type_cast_586_inst_req_1 : boolean;
  signal type_cast_599_inst_req_0 : boolean;
  signal type_cast_658_inst_ack_1 : boolean;
  signal type_cast_574_inst_ack_1 : boolean;
  signal type_cast_524_inst_ack_0 : boolean;
  signal type_cast_536_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_req_0 : boolean;
  signal type_cast_549_inst_ack_1 : boolean;
  signal type_cast_658_inst_ack_0 : boolean;
  signal type_cast_1103_inst_ack_0 : boolean;
  signal type_cast_611_inst_ack_0 : boolean;
  signal type_cast_599_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_545_inst_ack_0 : boolean;
  signal type_cast_636_inst_req_1 : boolean;
  signal type_cast_549_inst_req_0 : boolean;
  signal type_cast_536_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_620_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_620_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_595_inst_req_0 : boolean;
  signal type_cast_524_inst_req_1 : boolean;
  signal type_cast_1205_inst_ack_0 : boolean;
  signal if_stmt_686_branch_ack_1 : boolean;
  signal type_cast_1005_inst_ack_0 : boolean;
  signal if_stmt_1053_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1298_inst_ack_1 : boolean;
  signal array_obj_ref_1092_index_offset_ack_1 : boolean;
  signal type_cast_678_inst_req_1 : boolean;
  signal ptr_deref_1096_store_0_req_0 : boolean;
  signal type_cast_662_inst_ack_1 : boolean;
  signal type_cast_1320_inst_ack_0 : boolean;
  signal type_cast_636_inst_ack_1 : boolean;
  signal if_stmt_686_branch_req_0 : boolean;
  signal type_cast_1302_inst_req_1 : boolean;
  signal array_obj_ref_1245_index_offset_req_0 : boolean;
  signal type_cast_1302_inst_req_0 : boolean;
  signal type_cast_1302_inst_ack_0 : boolean;
  signal if_stmt_686_branch_ack_0 : boolean;
  signal type_cast_706_inst_req_0 : boolean;
  signal type_cast_706_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1298_inst_req_1 : boolean;
  signal type_cast_706_inst_req_1 : boolean;
  signal type_cast_706_inst_ack_1 : boolean;
  signal type_cast_1174_inst_ack_0 : boolean;
  signal type_cast_574_inst_req_0 : boolean;
  signal type_cast_678_inst_req_0 : boolean;
  signal type_cast_1174_inst_req_0 : boolean;
  signal type_cast_624_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_ack_1 : boolean;
  signal type_cast_678_inst_ack_1 : boolean;
  signal type_cast_662_inst_ack_0 : boolean;
  signal type_cast_1103_inst_req_0 : boolean;
  signal type_cast_1205_inst_req_0 : boolean;
  signal type_cast_662_inst_req_0 : boolean;
  signal type_cast_649_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_595_inst_ack_1 : boolean;
  signal type_cast_649_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_645_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_645_inst_req_0 : boolean;
  signal array_obj_ref_1245_index_offset_ack_0 : boolean;
  signal type_cast_624_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_595_inst_req_1 : boolean;
  signal type_cast_611_inst_ack_1 : boolean;
  signal type_cast_511_inst_ack_1 : boolean;
  signal type_cast_611_inst_req_1 : boolean;
  signal type_cast_524_inst_ack_1 : boolean;
  signal type_cast_1046_inst_req_0 : boolean;
  signal type_cast_1103_inst_req_1 : boolean;
  signal if_stmt_1053_branch_ack_0 : boolean;
  signal type_cast_1174_inst_req_1 : boolean;
  signal type_cast_1103_inst_ack_1 : boolean;
  signal type_cast_1046_inst_ack_0 : boolean;
  signal addr_of_1246_final_reg_req_0 : boolean;
  signal array_obj_ref_1245_index_offset_req_1 : boolean;
  signal addr_of_1093_final_reg_req_0 : boolean;
  signal addr_of_1093_final_reg_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_457_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_457_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_457_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_457_inst_ack_1 : boolean;
  signal type_cast_461_inst_req_0 : boolean;
  signal type_cast_461_inst_ack_0 : boolean;
  signal type_cast_461_inst_req_1 : boolean;
  signal type_cast_461_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_470_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_470_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_470_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_470_inst_ack_1 : boolean;
  signal type_cast_474_inst_req_0 : boolean;
  signal type_cast_474_inst_ack_0 : boolean;
  signal type_cast_474_inst_req_1 : boolean;
  signal type_cast_474_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_482_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_482_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_482_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_482_inst_ack_1 : boolean;
  signal type_cast_486_inst_req_0 : boolean;
  signal type_cast_486_inst_ack_0 : boolean;
  signal type_cast_486_inst_req_1 : boolean;
  signal type_cast_486_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_495_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_495_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_495_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_495_inst_ack_1 : boolean;
  signal type_cast_499_inst_req_0 : boolean;
  signal type_cast_499_inst_ack_0 : boolean;
  signal type_cast_499_inst_req_1 : boolean;
  signal type_cast_499_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_507_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_507_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_507_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_507_inst_ack_1 : boolean;
  signal type_cast_511_inst_req_0 : boolean;
  signal type_cast_511_inst_ack_0 : boolean;
  signal type_cast_511_inst_req_1 : boolean;
  signal type_cast_722_inst_req_0 : boolean;
  signal type_cast_722_inst_ack_0 : boolean;
  signal type_cast_722_inst_req_1 : boolean;
  signal type_cast_722_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_req_0 : boolean;
  signal type_cast_731_inst_req_0 : boolean;
  signal type_cast_731_inst_ack_0 : boolean;
  signal type_cast_731_inst_req_1 : boolean;
  signal type_cast_731_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1316_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1298_inst_ack_0 : boolean;
  signal type_cast_1196_inst_ack_1 : boolean;
  signal type_cast_1196_inst_req_1 : boolean;
  signal type_cast_1253_inst_ack_1 : boolean;
  signal if_stmt_1153_branch_ack_0 : boolean;
  signal type_cast_1253_inst_req_1 : boolean;
  signal type_cast_741_inst_req_0 : boolean;
  signal type_cast_741_inst_ack_0 : boolean;
  signal type_cast_741_inst_req_1 : boolean;
  signal type_cast_741_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1316_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1298_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_ack_1 : boolean;
  signal array_obj_ref_1245_index_offset_ack_1 : boolean;
  signal type_cast_1196_inst_ack_0 : boolean;
  signal type_cast_1196_inst_req_0 : boolean;
  signal array_obj_ref_776_index_offset_req_0 : boolean;
  signal if_stmt_1153_branch_ack_1 : boolean;
  signal array_obj_ref_776_index_offset_ack_0 : boolean;
  signal array_obj_ref_776_index_offset_req_1 : boolean;
  signal array_obj_ref_776_index_offset_ack_1 : boolean;
  signal phi_stmt_1006_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_req_1 : boolean;
  signal if_stmt_1153_branch_req_0 : boolean;
  signal addr_of_777_final_reg_req_0 : boolean;
  signal addr_of_777_final_reg_ack_0 : boolean;
  signal type_cast_1253_inst_ack_0 : boolean;
  signal addr_of_777_final_reg_req_1 : boolean;
  signal addr_of_777_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_780_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_780_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_780_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_780_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_ack_0 : boolean;
  signal type_cast_1253_inst_req_0 : boolean;
  signal type_cast_784_inst_req_0 : boolean;
  signal type_cast_784_inst_ack_0 : boolean;
  signal type_cast_784_inst_req_1 : boolean;
  signal type_cast_784_inst_ack_1 : boolean;
  signal type_cast_1005_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_793_inst_req_0 : boolean;
  signal type_cast_1115_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_793_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_793_inst_req_1 : boolean;
  signal type_cast_1115_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_793_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_req_0 : boolean;
  signal type_cast_797_inst_req_0 : boolean;
  signal type_cast_797_inst_ack_0 : boolean;
  signal type_cast_797_inst_req_1 : boolean;
  signal type_cast_797_inst_ack_1 : boolean;
  signal type_cast_1187_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_811_inst_req_0 : boolean;
  signal type_cast_1115_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_811_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_811_inst_req_1 : boolean;
  signal type_cast_1115_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_811_inst_ack_1 : boolean;
  signal type_cast_1187_inst_req_1 : boolean;
  signal type_cast_815_inst_req_0 : boolean;
  signal type_cast_815_inst_ack_0 : boolean;
  signal type_cast_815_inst_req_1 : boolean;
  signal type_cast_815_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_829_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_829_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_829_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_829_inst_ack_1 : boolean;
  signal type_cast_1266_inst_ack_1 : boolean;
  signal type_cast_1187_inst_ack_0 : boolean;
  signal type_cast_1187_inst_req_0 : boolean;
  signal type_cast_1266_inst_req_1 : boolean;
  signal type_cast_833_inst_req_0 : boolean;
  signal type_cast_833_inst_ack_0 : boolean;
  signal type_cast_833_inst_req_1 : boolean;
  signal type_cast_833_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1316_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_req_1 : boolean;
  signal type_cast_1111_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_ack_1 : boolean;
  signal type_cast_1005_inst_req_1 : boolean;
  signal type_cast_1266_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1249_inst_ack_1 : boolean;
  signal type_cast_851_inst_req_0 : boolean;
  signal type_cast_1111_inst_req_1 : boolean;
  signal type_cast_851_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1249_inst_req_1 : boolean;
  signal type_cast_851_inst_req_1 : boolean;
  signal type_cast_851_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1316_inst_req_0 : boolean;
  signal type_cast_1210_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_865_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_865_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_865_inst_req_1 : boolean;
  signal type_cast_1111_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_865_inst_ack_1 : boolean;
  signal type_cast_1266_inst_req_0 : boolean;
  signal type_cast_869_inst_req_0 : boolean;
  signal type_cast_1111_inst_req_0 : boolean;
  signal type_cast_869_inst_ack_0 : boolean;
  signal type_cast_869_inst_req_1 : boolean;
  signal type_cast_869_inst_ack_1 : boolean;
  signal type_cast_1320_inst_ack_1 : boolean;
  signal type_cast_1284_inst_ack_1 : boolean;
  signal type_cast_1210_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_883_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_883_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_883_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_883_inst_ack_1 : boolean;
  signal type_cast_1178_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1249_inst_ack_0 : boolean;
  signal type_cast_887_inst_req_0 : boolean;
  signal type_cast_887_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1249_inst_req_0 : boolean;
  signal type_cast_887_inst_req_1 : boolean;
  signal type_cast_887_inst_ack_1 : boolean;
  signal type_cast_1284_inst_req_1 : boolean;
  signal type_cast_1320_inst_req_1 : boolean;
  signal type_cast_1178_inst_req_1 : boolean;
  signal type_cast_1210_inst_ack_0 : boolean;
  signal type_cast_1210_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_901_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_901_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_901_inst_req_1 : boolean;
  signal type_cast_1107_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_901_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1262_inst_ack_1 : boolean;
  signal type_cast_905_inst_req_0 : boolean;
  signal type_cast_1107_inst_req_1 : boolean;
  signal type_cast_905_inst_ack_0 : boolean;
  signal type_cast_905_inst_req_1 : boolean;
  signal type_cast_905_inst_ack_1 : boolean;
  signal type_cast_1284_inst_ack_0 : boolean;
  signal type_cast_1178_inst_ack_0 : boolean;
  signal type_cast_1178_inst_req_0 : boolean;
  signal type_cast_1107_inst_ack_0 : boolean;
  signal type_cast_1302_inst_ack_1 : boolean;
  signal array_obj_ref_1092_index_offset_req_1 : boolean;
  signal type_cast_1107_inst_req_0 : boolean;
  signal ptr_deref_913_store_0_req_0 : boolean;
  signal ptr_deref_913_store_0_ack_0 : boolean;
  signal if_stmt_1053_branch_req_0 : boolean;
  signal ptr_deref_913_store_0_req_1 : boolean;
  signal ptr_deref_913_store_0_ack_1 : boolean;
  signal type_cast_1284_inst_req_0 : boolean;
  signal type_cast_1320_inst_req_0 : boolean;
  signal addr_of_1093_final_reg_ack_1 : boolean;
  signal addr_of_1093_final_reg_req_1 : boolean;
  signal if_stmt_927_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1262_inst_req_1 : boolean;
  signal if_stmt_927_branch_ack_1 : boolean;
  signal ptr_deref_1096_store_0_ack_1 : boolean;
  signal if_stmt_927_branch_ack_0 : boolean;
  signal type_cast_1174_inst_ack_1 : boolean;
  signal array_obj_ref_1092_index_offset_ack_0 : boolean;
  signal type_cast_1046_inst_ack_1 : boolean;
  signal ptr_deref_1096_store_0_req_1 : boolean;
  signal addr_of_1246_final_reg_ack_1 : boolean;
  signal if_stmt_978_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1262_inst_ack_0 : boolean;
  signal type_cast_1046_inst_req_1 : boolean;
  signal if_stmt_978_branch_ack_1 : boolean;
  signal if_stmt_978_branch_ack_0 : boolean;
  signal addr_of_1246_final_reg_ack_0 : boolean;
  signal array_obj_ref_1092_index_offset_req_0 : boolean;
  signal type_cast_1205_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1262_inst_req_0 : boolean;
  signal addr_of_1246_final_reg_req_1 : boolean;
  signal type_cast_1205_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1027_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1027_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1027_inst_req_1 : boolean;
  signal type_cast_1005_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1027_inst_ack_1 : boolean;
  signal phi_stmt_958_req_1 : boolean;
  signal phi_stmt_999_req_1 : boolean;
  signal type_cast_1031_inst_req_0 : boolean;
  signal type_cast_1031_inst_ack_0 : boolean;
  signal type_cast_1031_inst_req_1 : boolean;
  signal type_cast_1031_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_ack_1 : boolean;
  signal phi_stmt_764_ack_0 : boolean;
  signal phi_stmt_764_req_0 : boolean;
  signal type_cast_767_inst_ack_1 : boolean;
  signal type_cast_1338_inst_req_0 : boolean;
  signal type_cast_1338_inst_ack_0 : boolean;
  signal phi_stmt_1427_req_1 : boolean;
  signal type_cast_1338_inst_req_1 : boolean;
  signal type_cast_1338_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1352_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1352_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1352_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1352_inst_ack_1 : boolean;
  signal type_cast_1239_inst_ack_0 : boolean;
  signal type_cast_1239_inst_req_0 : boolean;
  signal type_cast_1356_inst_req_0 : boolean;
  signal type_cast_1356_inst_ack_0 : boolean;
  signal type_cast_1356_inst_req_1 : boolean;
  signal type_cast_1356_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1370_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1370_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1370_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1370_inst_ack_1 : boolean;
  signal phi_stmt_1479_req_0 : boolean;
  signal type_cast_1374_inst_req_0 : boolean;
  signal type_cast_1374_inst_ack_0 : boolean;
  signal type_cast_1374_inst_req_1 : boolean;
  signal phi_stmt_1060_ack_0 : boolean;
  signal type_cast_1374_inst_ack_1 : boolean;
  signal phi_stmt_1006_req_0 : boolean;
  signal type_cast_1012_inst_ack_1 : boolean;
  signal phi_stmt_1060_req_0 : boolean;
  signal type_cast_1063_inst_ack_1 : boolean;
  signal ptr_deref_1382_store_0_req_0 : boolean;
  signal ptr_deref_1382_store_0_ack_0 : boolean;
  signal type_cast_767_inst_req_1 : boolean;
  signal ptr_deref_1382_store_0_req_1 : boolean;
  signal ptr_deref_1382_store_0_ack_1 : boolean;
  signal phi_stmt_1472_req_1 : boolean;
  signal type_cast_1478_inst_ack_1 : boolean;
  signal type_cast_1012_inst_req_1 : boolean;
  signal if_stmt_1396_branch_req_0 : boolean;
  signal type_cast_767_inst_ack_0 : boolean;
  signal if_stmt_1396_branch_ack_1 : boolean;
  signal type_cast_767_inst_req_0 : boolean;
  signal if_stmt_1396_branch_ack_0 : boolean;
  signal type_cast_1012_inst_ack_0 : boolean;
  signal phi_stmt_1472_req_0 : boolean;
  signal type_cast_1012_inst_req_0 : boolean;
  signal phi_stmt_1427_req_0 : boolean;
  signal if_stmt_1447_branch_req_0 : boolean;
  signal phi_stmt_999_req_0 : boolean;
  signal if_stmt_1447_branch_ack_1 : boolean;
  signal if_stmt_1447_branch_ack_0 : boolean;
  signal phi_stmt_1233_ack_0 : boolean;
  signal type_cast_1430_inst_ack_1 : boolean;
  signal type_cast_1462_inst_req_0 : boolean;
  signal type_cast_1063_inst_req_1 : boolean;
  signal type_cast_1462_inst_ack_0 : boolean;
  signal type_cast_1430_inst_req_1 : boolean;
  signal type_cast_1462_inst_req_1 : boolean;
  signal type_cast_1462_inst_ack_1 : boolean;
  signal type_cast_1478_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1500_inst_req_0 : boolean;
  signal type_cast_1063_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1500_inst_ack_0 : boolean;
  signal phi_stmt_1233_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1500_inst_req_1 : boolean;
  signal type_cast_1063_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1500_inst_ack_1 : boolean;
  signal type_cast_1504_inst_req_0 : boolean;
  signal type_cast_1504_inst_ack_0 : boolean;
  signal phi_stmt_1233_req_1 : boolean;
  signal type_cast_1504_inst_req_1 : boolean;
  signal type_cast_1504_inst_ack_1 : boolean;
  signal type_cast_1478_inst_ack_0 : boolean;
  signal type_cast_1430_inst_ack_0 : boolean;
  signal type_cast_1519_inst_req_0 : boolean;
  signal type_cast_1519_inst_ack_0 : boolean;
  signal type_cast_1430_inst_req_0 : boolean;
  signal type_cast_1519_inst_req_1 : boolean;
  signal type_cast_1519_inst_ack_1 : boolean;
  signal type_cast_1478_inst_req_0 : boolean;
  signal if_stmt_1526_branch_req_0 : boolean;
  signal if_stmt_1526_branch_ack_1 : boolean;
  signal if_stmt_1526_branch_ack_0 : boolean;
  signal phi_stmt_764_req_1 : boolean;
  signal type_cast_1239_inst_ack_1 : boolean;
  signal array_obj_ref_1565_index_offset_req_0 : boolean;
  signal array_obj_ref_1565_index_offset_ack_0 : boolean;
  signal array_obj_ref_1565_index_offset_req_1 : boolean;
  signal array_obj_ref_1565_index_offset_ack_1 : boolean;
  signal addr_of_1566_final_reg_req_0 : boolean;
  signal addr_of_1566_final_reg_ack_0 : boolean;
  signal addr_of_1566_final_reg_req_1 : boolean;
  signal addr_of_1566_final_reg_ack_1 : boolean;
  signal phi_stmt_958_ack_0 : boolean;
  signal phi_stmt_958_req_0 : boolean;
  signal type_cast_961_inst_ack_1 : boolean;
  signal type_cast_961_inst_req_1 : boolean;
  signal type_cast_961_inst_ack_0 : boolean;
  signal type_cast_961_inst_req_0 : boolean;
  signal ptr_deref_1569_store_0_req_0 : boolean;
  signal ptr_deref_1569_store_0_ack_0 : boolean;
  signal ptr_deref_1569_store_0_req_1 : boolean;
  signal ptr_deref_1569_store_0_ack_1 : boolean;
  signal phi_stmt_1006_ack_0 : boolean;
  signal type_cast_1239_inst_req_1 : boolean;
  signal phi_stmt_999_ack_0 : boolean;
  signal call_stmt_1576_call_req_0 : boolean;
  signal call_stmt_1576_call_ack_0 : boolean;
  signal call_stmt_1576_call_req_1 : boolean;
  signal call_stmt_1576_call_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1583_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1583_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1583_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1583_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1587_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1587_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1587_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1587_inst_ack_1 : boolean;
  signal type_cast_1616_inst_req_0 : boolean;
  signal type_cast_1616_inst_ack_0 : boolean;
  signal type_cast_1616_inst_req_1 : boolean;
  signal type_cast_1616_inst_ack_1 : boolean;
  signal type_cast_1626_inst_req_0 : boolean;
  signal type_cast_1626_inst_ack_0 : boolean;
  signal type_cast_1626_inst_req_1 : boolean;
  signal type_cast_1626_inst_ack_1 : boolean;
  signal type_cast_1635_inst_req_0 : boolean;
  signal type_cast_1635_inst_ack_0 : boolean;
  signal type_cast_1635_inst_req_1 : boolean;
  signal type_cast_1635_inst_ack_1 : boolean;
  signal type_cast_1664_inst_req_0 : boolean;
  signal type_cast_1664_inst_ack_0 : boolean;
  signal type_cast_1664_inst_req_1 : boolean;
  signal type_cast_1664_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1666_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_1666_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1666_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_1666_inst_ack_1 : boolean;
  signal type_cast_1671_inst_req_0 : boolean;
  signal type_cast_1671_inst_ack_0 : boolean;
  signal type_cast_1671_inst_req_1 : boolean;
  signal type_cast_1671_inst_ack_1 : boolean;
  signal type_cast_1675_inst_req_0 : boolean;
  signal type_cast_1675_inst_ack_0 : boolean;
  signal type_cast_1675_inst_req_1 : boolean;
  signal type_cast_1675_inst_ack_1 : boolean;
  signal call_stmt_1686_call_req_0 : boolean;
  signal call_stmt_1686_call_ack_0 : boolean;
  signal call_stmt_1686_call_req_1 : boolean;
  signal call_stmt_1686_call_ack_1 : boolean;
  signal call_stmt_1693_call_req_0 : boolean;
  signal call_stmt_1693_call_ack_0 : boolean;
  signal call_stmt_1693_call_req_1 : boolean;
  signal call_stmt_1693_call_ack_1 : boolean;
  signal if_stmt_1705_branch_req_0 : boolean;
  signal if_stmt_1705_branch_ack_1 : boolean;
  signal if_stmt_1705_branch_ack_0 : boolean;
  signal type_cast_1715_inst_req_0 : boolean;
  signal type_cast_1715_inst_ack_0 : boolean;
  signal type_cast_1715_inst_req_1 : boolean;
  signal type_cast_1715_inst_ack_1 : boolean;
  signal call_stmt_1719_call_req_0 : boolean;
  signal call_stmt_1719_call_ack_0 : boolean;
  signal call_stmt_1719_call_req_1 : boolean;
  signal call_stmt_1719_call_ack_1 : boolean;
  signal type_cast_1723_inst_req_0 : boolean;
  signal type_cast_1723_inst_ack_0 : boolean;
  signal type_cast_1723_inst_req_1 : boolean;
  signal type_cast_1723_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1730_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1730_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1730_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1730_inst_ack_1 : boolean;
  signal type_cast_1485_inst_req_0 : boolean;
  signal type_cast_1485_inst_ack_0 : boolean;
  signal type_cast_1485_inst_req_1 : boolean;
  signal type_cast_1485_inst_ack_1 : boolean;
  signal phi_stmt_1479_req_1 : boolean;
  signal phi_stmt_1472_ack_0 : boolean;
  signal phi_stmt_1479_ack_0 : boolean;
  signal type_cast_1536_inst_req_0 : boolean;
  signal type_cast_1536_inst_ack_0 : boolean;
  signal type_cast_1536_inst_req_1 : boolean;
  signal type_cast_1536_inst_ack_1 : boolean;
  signal phi_stmt_1533_req_0 : boolean;
  signal phi_stmt_1533_ack_0 : boolean;
  signal phi_stmt_1644_req_1 : boolean;
  signal type_cast_1647_inst_req_0 : boolean;
  signal type_cast_1647_inst_ack_0 : boolean;
  signal type_cast_1647_inst_req_1 : boolean;
  signal type_cast_1647_inst_ack_1 : boolean;
  signal phi_stmt_1644_req_0 : boolean;
  signal phi_stmt_1644_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_1129_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1129_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_1129_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1129_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_1129: Block -- control-path 
    signal convolution3D_CP_1129_elements: BooleanArray(337 downto 0);
    -- 
  begin -- 
    convolution3D_CP_1129_elements(0) <= convolution3D_CP_1129_start;
    convolution3D_CP_1129_symbol <= convolution3D_CP_1129_elements(269);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	73 
    -- CP-element group 0:  members (65) 
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_454/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/branch_block_stmt_454__entry__
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685__entry__
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_update_start_
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_Update/cr
      -- 
    cr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_649_inst_req_1); -- 
    cr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_536_inst_req_1); -- 
    cr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_574_inst_req_1); -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_561_inst_req_1); -- 
    cr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_549_inst_req_1); -- 
    cr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_658_inst_req_1); -- 
    cr_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_662_inst_req_1); -- 
    cr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_586_inst_req_1); -- 
    cr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_599_inst_req_1); -- 
    cr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_636_inst_req_1); -- 
    cr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_524_inst_req_1); -- 
    cr_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_678_inst_req_1); -- 
    cr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_624_inst_req_1); -- 
    cr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_611_inst_req_1); -- 
    rr_1245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => RPIPE_maxpool_input_pipe_457_inst_req_0); -- 
    cr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_461_inst_req_1); -- 
    cr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_474_inst_req_1); -- 
    cr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_486_inst_req_1); -- 
    cr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_499_inst_req_1); -- 
    cr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_511_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_update_start_
      -- CP-element group 1: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_Update/cr
      -- 
    ra_1246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_457_inst_ack_0, ack => convolution3D_CP_1129_elements(1)); -- 
    cr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(1), ack => RPIPE_maxpool_input_pipe_457_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_457_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_Sample/rr
      -- 
    ca_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_457_inst_ack_1, ack => convolution3D_CP_1129_elements(2)); -- 
    rr_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(2), ack => type_cast_461_inst_req_0); -- 
    rr_1273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(2), ack => RPIPE_maxpool_input_pipe_470_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_Sample/ra
      -- 
    ra_1260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_0, ack => convolution3D_CP_1129_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_461_Update/ca
      -- 
    ca_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_1, ack => convolution3D_CP_1129_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_update_start_
      -- CP-element group 5: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_Update/cr
      -- 
    ra_1274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_470_inst_ack_0, ack => convolution3D_CP_1129_elements(5)); -- 
    cr_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(5), ack => RPIPE_maxpool_input_pipe_470_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_470_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_Sample/rr
      -- 
    ca_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_470_inst_ack_1, ack => convolution3D_CP_1129_elements(6)); -- 
    rr_1287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(6), ack => type_cast_474_inst_req_0); -- 
    rr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(6), ack => RPIPE_maxpool_input_pipe_482_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_Sample/ra
      -- 
    ra_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_474_inst_ack_0, ack => convolution3D_CP_1129_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_474_Update/ca
      -- 
    ca_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_474_inst_ack_1, ack => convolution3D_CP_1129_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_update_start_
      -- CP-element group 9: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_Update/cr
      -- 
    ra_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_482_inst_ack_0, ack => convolution3D_CP_1129_elements(9)); -- 
    cr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(9), ack => RPIPE_maxpool_input_pipe_482_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_482_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_Sample/rr
      -- 
    ca_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_482_inst_ack_1, ack => convolution3D_CP_1129_elements(10)); -- 
    rr_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(10), ack => type_cast_486_inst_req_0); -- 
    rr_1329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(10), ack => RPIPE_maxpool_input_pipe_495_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_Sample/ra
      -- 
    ra_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_0, ack => convolution3D_CP_1129_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_486_Update/ca
      -- 
    ca_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_1, ack => convolution3D_CP_1129_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_update_start_
      -- CP-element group 13: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_Update/cr
      -- 
    ra_1330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_495_inst_ack_0, ack => convolution3D_CP_1129_elements(13)); -- 
    cr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(13), ack => RPIPE_maxpool_input_pipe_495_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_495_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_Sample/rr
      -- 
    ca_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_495_inst_ack_1, ack => convolution3D_CP_1129_elements(14)); -- 
    rr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(14), ack => type_cast_499_inst_req_0); -- 
    rr_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(14), ack => RPIPE_maxpool_input_pipe_507_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_Sample/ra
      -- 
    ra_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_499_inst_ack_0, ack => convolution3D_CP_1129_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_499_Update/ca
      -- 
    ca_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_499_inst_ack_1, ack => convolution3D_CP_1129_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_update_start_
      -- CP-element group 17: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_Update/cr
      -- 
    ra_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_507_inst_ack_0, ack => convolution3D_CP_1129_elements(17)); -- 
    cr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(17), ack => RPIPE_maxpool_input_pipe_507_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_507_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_Sample/rr
      -- 
    ca_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_507_inst_ack_1, ack => convolution3D_CP_1129_elements(18)); -- 
    rr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(18), ack => type_cast_511_inst_req_0); -- 
    rr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(18), ack => RPIPE_maxpool_input_pipe_520_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_Sample/ra
      -- 
    ra_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_511_inst_ack_0, ack => convolution3D_CP_1129_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_511_Update/$exit
      -- 
    ca_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_511_inst_ack_1, ack => convolution3D_CP_1129_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_update_start_
      -- CP-element group 21: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_sample_completed_
      -- 
    ra_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_520_inst_ack_0, ack => convolution3D_CP_1129_elements(21)); -- 
    cr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(21), ack => RPIPE_maxpool_input_pipe_520_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_520_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_sample_start_
      -- 
    ca_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_520_inst_ack_1, ack => convolution3D_CP_1129_elements(22)); -- 
    rr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(22), ack => type_cast_524_inst_req_0); -- 
    rr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(22), ack => RPIPE_maxpool_input_pipe_532_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_Sample/ra
      -- 
    ra_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_524_inst_ack_0, ack => convolution3D_CP_1129_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_524_Update/ca
      -- 
    ca_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_524_inst_ack_1, ack => convolution3D_CP_1129_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_update_start_
      -- CP-element group 25: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_sample_completed_
      -- 
    ra_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_532_inst_ack_0, ack => convolution3D_CP_1129_elements(25)); -- 
    cr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(25), ack => RPIPE_maxpool_input_pipe_532_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_532_update_completed_
      -- 
    ca_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_532_inst_ack_1, ack => convolution3D_CP_1129_elements(26)); -- 
    rr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(26), ack => type_cast_536_inst_req_0); -- 
    rr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(26), ack => RPIPE_maxpool_input_pipe_545_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_sample_completed_
      -- 
    ra_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_536_inst_ack_0, ack => convolution3D_CP_1129_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	74 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_536_update_completed_
      -- 
    ca_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_536_inst_ack_1, ack => convolution3D_CP_1129_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_Update/cr
      -- CP-element group 29: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_update_start_
      -- 
    ra_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_545_inst_ack_0, ack => convolution3D_CP_1129_elements(29)); -- 
    cr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(29), ack => RPIPE_maxpool_input_pipe_545_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_545_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_Sample/$entry
      -- 
    ca_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_545_inst_ack_1, ack => convolution3D_CP_1129_elements(30)); -- 
    rr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(30), ack => type_cast_549_inst_req_0); -- 
    rr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(30), ack => RPIPE_maxpool_input_pipe_557_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_sample_completed_
      -- 
    ra_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_549_inst_ack_0, ack => convolution3D_CP_1129_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	74 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_549_update_completed_
      -- 
    ca_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_549_inst_ack_1, ack => convolution3D_CP_1129_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_update_start_
      -- CP-element group 33: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_Update/$entry
      -- 
    ra_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_557_inst_ack_0, ack => convolution3D_CP_1129_elements(33)); -- 
    cr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(33), ack => RPIPE_maxpool_input_pipe_557_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_557_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_sample_start_
      -- 
    ca_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_557_inst_ack_1, ack => convolution3D_CP_1129_elements(34)); -- 
    rr_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(34), ack => type_cast_561_inst_req_0); -- 
    rr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(34), ack => RPIPE_maxpool_input_pipe_570_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_sample_completed_
      -- 
    ra_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_0, ack => convolution3D_CP_1129_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	74 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_561_update_completed_
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_1, ack => convolution3D_CP_1129_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_update_start_
      -- CP-element group 37: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_sample_completed_
      -- 
    ra_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_570_inst_ack_0, ack => convolution3D_CP_1129_elements(37)); -- 
    cr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(37), ack => RPIPE_maxpool_input_pipe_570_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_570_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_Sample/rr
      -- 
    ca_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_570_inst_ack_1, ack => convolution3D_CP_1129_elements(38)); -- 
    rr_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(38), ack => type_cast_574_inst_req_0); -- 
    rr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(38), ack => RPIPE_maxpool_input_pipe_582_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_Sample/$exit
      -- 
    ra_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_0, ack => convolution3D_CP_1129_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	74 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_574_update_completed_
      -- 
    ca_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_1, ack => convolution3D_CP_1129_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_update_start_
      -- CP-element group 41: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_Update/$entry
      -- 
    ra_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_582_inst_ack_0, ack => convolution3D_CP_1129_elements(41)); -- 
    cr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(41), ack => RPIPE_maxpool_input_pipe_582_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_582_Update/ca
      -- 
    ca_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_582_inst_ack_1, ack => convolution3D_CP_1129_elements(42)); -- 
    rr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(42), ack => type_cast_586_inst_req_0); -- 
    rr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(42), ack => RPIPE_maxpool_input_pipe_595_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_sample_completed_
      -- 
    ra_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_586_inst_ack_0, ack => convolution3D_CP_1129_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	74 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_586_update_completed_
      -- 
    ca_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_586_inst_ack_1, ack => convolution3D_CP_1129_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_update_start_
      -- CP-element group 45: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_Update/cr
      -- 
    ra_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_595_inst_ack_0, ack => convolution3D_CP_1129_elements(45)); -- 
    cr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(45), ack => RPIPE_maxpool_input_pipe_595_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_595_Update/ca
      -- 
    ca_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_595_inst_ack_1, ack => convolution3D_CP_1129_elements(46)); -- 
    rr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(46), ack => type_cast_599_inst_req_0); -- 
    rr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(46), ack => RPIPE_maxpool_input_pipe_607_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_sample_completed_
      -- 
    ra_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_599_inst_ack_0, ack => convolution3D_CP_1129_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_599_Update/$exit
      -- 
    ca_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_599_inst_ack_1, ack => convolution3D_CP_1129_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_update_start_
      -- CP-element group 49: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_Update/cr
      -- 
    ra_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_607_inst_ack_0, ack => convolution3D_CP_1129_elements(49)); -- 
    cr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(49), ack => RPIPE_maxpool_input_pipe_607_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_607_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_sample_start_
      -- 
    ca_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_607_inst_ack_1, ack => convolution3D_CP_1129_elements(50)); -- 
    rr_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(50), ack => type_cast_611_inst_req_0); -- 
    rr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(50), ack => RPIPE_maxpool_input_pipe_620_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_sample_completed_
      -- 
    ra_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_611_inst_ack_0, ack => convolution3D_CP_1129_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	74 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_611_Update/ca
      -- 
    ca_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_611_inst_ack_1, ack => convolution3D_CP_1129_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_update_start_
      -- CP-element group 53: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_Update/cr
      -- 
    ra_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_620_inst_ack_0, ack => convolution3D_CP_1129_elements(53)); -- 
    cr_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(53), ack => RPIPE_maxpool_input_pipe_620_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_620_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_sample_start_
      -- 
    ca_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_620_inst_ack_1, ack => convolution3D_CP_1129_elements(54)); -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(54), ack => type_cast_624_inst_req_0); -- 
    rr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(54), ack => RPIPE_maxpool_input_pipe_632_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_sample_completed_
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_624_inst_ack_0, ack => convolution3D_CP_1129_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	74 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_624_Update/$exit
      -- 
    ca_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_624_inst_ack_1, ack => convolution3D_CP_1129_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_update_start_
      -- CP-element group 57: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_sample_completed_
      -- 
    ra_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_632_inst_ack_0, ack => convolution3D_CP_1129_elements(57)); -- 
    cr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(57), ack => RPIPE_maxpool_input_pipe_632_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_632_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_Sample/rr
      -- 
    ca_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_632_inst_ack_1, ack => convolution3D_CP_1129_elements(58)); -- 
    rr_1651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(58), ack => type_cast_636_inst_req_0); -- 
    rr_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(58), ack => RPIPE_maxpool_input_pipe_645_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_Sample/ra
      -- 
    ra_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_0, ack => convolution3D_CP_1129_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_636_Update/ca
      -- 
    ca_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_1, ack => convolution3D_CP_1129_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_Update/cr
      -- CP-element group 61: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_update_start_
      -- CP-element group 61: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_Sample/ra
      -- 
    ra_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_645_inst_ack_0, ack => convolution3D_CP_1129_elements(61)); -- 
    cr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(61), ack => RPIPE_maxpool_input_pipe_645_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/RPIPE_maxpool_input_pipe_645_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_Sample/rr
      -- 
    ca_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_645_inst_ack_1, ack => convolution3D_CP_1129_elements(62)); -- 
    rr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(62), ack => type_cast_649_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_Sample/ra
      -- 
    ra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_0, ack => convolution3D_CP_1129_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	74 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_649_update_completed_
      -- 
    ca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_1, ack => convolution3D_CP_1129_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	16 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_sample_start_
      -- 
    rr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(65), ack => type_cast_658_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(12) & convolution3D_CP_1129_elements(16);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_sample_completed_
      -- 
    ra_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_658_inst_ack_0, ack => convolution3D_CP_1129_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_658_update_completed_
      -- 
    ca_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_658_inst_ack_1, ack => convolution3D_CP_1129_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	20 
    -- CP-element group 68: 	24 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_Sample/rr
      -- 
    rr_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(68), ack => type_cast_662_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(20) & convolution3D_CP_1129_elements(24);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_Sample/ra
      -- 
    ra_1708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_662_inst_ack_0, ack => convolution3D_CP_1129_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_662_update_completed_
      -- 
    ca_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_662_inst_ack_1, ack => convolution3D_CP_1129_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	4 
    -- CP-element group 71: 	8 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_Sample/rr
      -- 
    rr_1721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(71), ack => type_cast_678_inst_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(4) & convolution3D_CP_1129_elements(8) & convolution3D_CP_1129_elements(67) & convolution3D_CP_1129_elements(70);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_Sample/$exit
      -- 
    ra_1722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_678_inst_ack_0, ack => convolution3D_CP_1129_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/type_cast_678_Update/ca
      -- 
    ca_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_678_inst_ack_1, ack => convolution3D_CP_1129_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: 	32 
    -- CP-element group 74: 	36 
    -- CP-element group 74: 	40 
    -- CP-element group 74: 	44 
    -- CP-element group 74: 	48 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	56 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	64 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_454/if_stmt_686_else_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_454/if_stmt_686_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_454/if_stmt_686_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_454/R_cmp325_687_place
      -- CP-element group 74: 	 branch_block_stmt_454/if_stmt_686_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_454/if_stmt_686_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_454/if_stmt_686_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685__exit__
      -- CP-element group 74: 	 branch_block_stmt_454/if_stmt_686__entry__
      -- CP-element group 74: 	 branch_block_stmt_454/assign_stmt_458_to_assign_stmt_685/$exit
      -- 
    branch_req_1735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(74), ack => if_stmt_686_branch_req_0); -- 
    convolution3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(28) & convolution3D_CP_1129_elements(32) & convolution3D_CP_1129_elements(36) & convolution3D_CP_1129_elements(40) & convolution3D_CP_1129_elements(44) & convolution3D_CP_1129_elements(48) & convolution3D_CP_1129_elements(52) & convolution3D_CP_1129_elements(56) & convolution3D_CP_1129_elements(60) & convolution3D_CP_1129_elements(64) & convolution3D_CP_1129_elements(73);
      gj_convolution3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	78 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	80 
    -- CP-element group 75: 	81 
    -- CP-element group 75: 	82 
    -- CP-element group 75: 	85 
    -- CP-element group 75:  members (33) 
      -- CP-element group 75: 	 branch_block_stmt_454/if_stmt_686_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_454/if_stmt_686_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_update_start_
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_454/entry_bbx_xnph327
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/$entry
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_update_start_
      -- CP-element group 75: 	 branch_block_stmt_454/merge_stmt_692__exit__
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761__entry__
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_update_start_
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_update_start_
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_454/entry_bbx_xnph327_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_454/entry_bbx_xnph327_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_454/merge_stmt_692_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_454/merge_stmt_692_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_454/merge_stmt_692_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_454/merge_stmt_692_PhiAck/dummy
      -- 
    if_choice_transition_1740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_686_branch_ack_1, ack => convolution3D_CP_1129_elements(75)); -- 
    rr_1757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_706_inst_req_0); -- 
    cr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_706_inst_req_1); -- 
    rr_1771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_722_inst_req_0); -- 
    cr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_722_inst_req_1); -- 
    rr_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_731_inst_req_0); -- 
    cr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_731_inst_req_1); -- 
    cr_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_741_inst_req_1); -- 
    -- CP-element group 76:  transition  place  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	276 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_454/entry_forx_xend
      -- CP-element group 76: 	 branch_block_stmt_454/if_stmt_686_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_454/if_stmt_686_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_454/entry_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_454/entry_forx_xend_PhiReq/phi_stmt_958/$entry
      -- CP-element group 76: 	 branch_block_stmt_454/entry_forx_xend_PhiReq/$entry
      -- 
    else_choice_transition_1744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_686_branch_ack_0, ack => convolution3D_CP_1129_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_sample_completed_
      -- 
    ra_1758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_706_inst_ack_0, ack => convolution3D_CP_1129_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	86 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_706_update_completed_
      -- 
    ca_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_706_inst_ack_1, ack => convolution3D_CP_1129_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_Sample/ra
      -- 
    ra_1772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_0, ack => convolution3D_CP_1129_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_722_Update/ca
      -- 
    ca_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_1, ack => convolution3D_CP_1129_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_Sample/ra
      -- 
    ra_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_0, ack => convolution3D_CP_1129_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	75 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_731_Update/ca
      -- 
    ca_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_1, ack => convolution3D_CP_1129_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_Sample/rr
      -- 
    rr_1799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(83), ack => type_cast_741_inst_req_0); -- 
    convolution3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(80) & convolution3D_CP_1129_elements(82);
      gj_convolution3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_Sample/ra
      -- 
    ra_1800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_741_inst_ack_0, ack => convolution3D_CP_1129_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	75 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/type_cast_741_Update/ca
      -- 
    ca_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_741_inst_ack_1, ack => convolution3D_CP_1129_elements(85)); -- 
    -- CP-element group 86:  join  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	78 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	270 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761/$exit
      -- CP-element group 86: 	 branch_block_stmt_454/assign_stmt_697_to_assign_stmt_761__exit__
      -- CP-element group 86: 	 branch_block_stmt_454/bbx_xnph327_forx_xbody
      -- CP-element group 86: 	 branch_block_stmt_454/bbx_xnph327_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_454/bbx_xnph327_forx_xbody_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_454/bbx_xnph327_forx_xbody_PhiReq/phi_stmt_764/$entry
      -- 
    convolution3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(78) & convolution3D_CP_1129_elements(85);
      gj_convolution3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	275 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	126 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_sample_complete
      -- CP-element group 87: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Sample/ack
      -- 
    ack_1834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_776_index_offset_ack_0, ack => convolution3D_CP_1129_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	275 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (11) 
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_offset_calculated
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_request/$entry
      -- CP-element group 88: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_request/req
      -- 
    ack_1839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_776_index_offset_ack_1, ack => convolution3D_CP_1129_elements(88)); -- 
    req_1848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(88), ack => addr_of_777_final_reg_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_request/$exit
      -- CP-element group 89: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_request/ack
      -- 
    ack_1849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_777_final_reg_ack_0, ack => convolution3D_CP_1129_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	275 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	123 
    -- CP-element group 90:  members (19) 
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_complete/ack
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_word_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_root_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_address_resized
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_addr_resize/$entry
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_addr_resize/$exit
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_addr_resize/base_resize_req
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_addr_resize/base_resize_ack
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_plus_offset/$entry
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_plus_offset/$exit
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_word_addrgen/$entry
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_word_addrgen/$exit
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_word_addrgen/root_register_req
      -- CP-element group 90: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_word_addrgen/root_register_ack
      -- 
    ack_1854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_777_final_reg_ack_1, ack => convolution3D_CP_1129_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	275 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_update_start_
      -- CP-element group 91: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_Update/cr
      -- 
    ra_1863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_780_inst_ack_0, ack => convolution3D_CP_1129_elements(91)); -- 
    cr_1867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(91), ack => RPIPE_maxpool_input_pipe_780_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_Sample/rr
      -- 
    ca_1868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_780_inst_ack_1, ack => convolution3D_CP_1129_elements(92)); -- 
    rr_1876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(92), ack => type_cast_784_inst_req_0); -- 
    rr_1890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(92), ack => RPIPE_maxpool_input_pipe_793_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_Sample/ra
      -- 
    ra_1877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_784_inst_ack_0, ack => convolution3D_CP_1129_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	275 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	123 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_Update/ca
      -- 
    ca_1882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_784_inst_ack_1, ack => convolution3D_CP_1129_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_update_start_
      -- CP-element group 95: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_Update/cr
      -- 
    ra_1891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_793_inst_ack_0, ack => convolution3D_CP_1129_elements(95)); -- 
    cr_1895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(95), ack => RPIPE_maxpool_input_pipe_793_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_793_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_Sample/rr
      -- 
    ca_1896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_793_inst_ack_1, ack => convolution3D_CP_1129_elements(96)); -- 
    rr_1904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(96), ack => type_cast_797_inst_req_0); -- 
    rr_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(96), ack => RPIPE_maxpool_input_pipe_811_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_Sample/ra
      -- 
    ra_1905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_797_inst_ack_0, ack => convolution3D_CP_1129_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	275 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	123 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_Update/ca
      -- 
    ca_1910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_797_inst_ack_1, ack => convolution3D_CP_1129_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_update_start_
      -- CP-element group 99: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_Update/cr
      -- 
    ra_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_811_inst_ack_0, ack => convolution3D_CP_1129_elements(99)); -- 
    cr_1923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(99), ack => RPIPE_maxpool_input_pipe_811_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_811_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_Sample/rr
      -- 
    ca_1924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_811_inst_ack_1, ack => convolution3D_CP_1129_elements(100)); -- 
    rr_1932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(100), ack => type_cast_815_inst_req_0); -- 
    rr_1946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(100), ack => RPIPE_maxpool_input_pipe_829_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_Sample/ra
      -- 
    ra_1933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_815_inst_ack_0, ack => convolution3D_CP_1129_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	275 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	123 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_Update/ca
      -- 
    ca_1938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_815_inst_ack_1, ack => convolution3D_CP_1129_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_update_start_
      -- CP-element group 103: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_Update/cr
      -- 
    ra_1947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_829_inst_ack_0, ack => convolution3D_CP_1129_elements(103)); -- 
    cr_1951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(103), ack => RPIPE_maxpool_input_pipe_829_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	107 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_829_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_Sample/rr
      -- 
    ca_1952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_829_inst_ack_1, ack => convolution3D_CP_1129_elements(104)); -- 
    rr_1960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(104), ack => type_cast_833_inst_req_0); -- 
    rr_1974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(104), ack => RPIPE_maxpool_input_pipe_847_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_Sample/ra
      -- 
    ra_1961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_0, ack => convolution3D_CP_1129_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	275 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	123 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_Update/ca
      -- 
    ca_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_1, ack => convolution3D_CP_1129_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_update_start_
      -- CP-element group 107: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_Update/cr
      -- 
    ra_1975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_847_inst_ack_0, ack => convolution3D_CP_1129_elements(107)); -- 
    cr_1979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(107), ack => RPIPE_maxpool_input_pipe_847_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_847_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_Sample/rr
      -- 
    ca_1980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_847_inst_ack_1, ack => convolution3D_CP_1129_elements(108)); -- 
    rr_1988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(108), ack => type_cast_851_inst_req_0); -- 
    rr_2002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(108), ack => RPIPE_maxpool_input_pipe_865_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_Sample/ra
      -- 
    ra_1989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_0, ack => convolution3D_CP_1129_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	275 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	123 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_Update/ca
      -- 
    ca_1994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_1, ack => convolution3D_CP_1129_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_update_start_
      -- CP-element group 111: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_Update/cr
      -- 
    ra_2003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_865_inst_ack_0, ack => convolution3D_CP_1129_elements(111)); -- 
    cr_2007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(111), ack => RPIPE_maxpool_input_pipe_865_inst_req_1); -- 
    -- CP-element group 112:  fork  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_865_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_Sample/rr
      -- 
    ca_2008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_865_inst_ack_1, ack => convolution3D_CP_1129_elements(112)); -- 
    rr_2016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(112), ack => type_cast_869_inst_req_0); -- 
    rr_2030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(112), ack => RPIPE_maxpool_input_pipe_883_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_Sample/ra
      -- 
    ra_2017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_869_inst_ack_0, ack => convolution3D_CP_1129_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	275 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	123 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_Update/ca
      -- 
    ca_2022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_869_inst_ack_1, ack => convolution3D_CP_1129_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_update_start_
      -- CP-element group 115: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_Update/cr
      -- 
    ra_2031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_883_inst_ack_0, ack => convolution3D_CP_1129_elements(115)); -- 
    cr_2035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(115), ack => RPIPE_maxpool_input_pipe_883_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_883_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_Sample/rr
      -- 
    ca_2036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_883_inst_ack_1, ack => convolution3D_CP_1129_elements(116)); -- 
    rr_2044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(116), ack => type_cast_887_inst_req_0); -- 
    rr_2058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(116), ack => RPIPE_maxpool_input_pipe_901_inst_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_Sample/ra
      -- 
    ra_2045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_0, ack => convolution3D_CP_1129_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	275 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_Update/ca
      -- 
    ca_2050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_1, ack => convolution3D_CP_1129_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_update_start_
      -- CP-element group 119: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_Update/cr
      -- 
    ra_2059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_901_inst_ack_0, ack => convolution3D_CP_1129_elements(119)); -- 
    cr_2063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(119), ack => RPIPE_maxpool_input_pipe_901_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_901_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_Sample/rr
      -- 
    ca_2064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_901_inst_ack_1, ack => convolution3D_CP_1129_elements(120)); -- 
    rr_2072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(120), ack => type_cast_905_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_Sample/ra
      -- 
    ra_2073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_0, ack => convolution3D_CP_1129_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	275 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_Update/ca
      -- 
    ca_2078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_1, ack => convolution3D_CP_1129_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	90 
    -- CP-element group 123: 	94 
    -- CP-element group 123: 	98 
    -- CP-element group 123: 	102 
    -- CP-element group 123: 	106 
    -- CP-element group 123: 	110 
    -- CP-element group 123: 	114 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (9) 
      -- CP-element group 123: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/ptr_deref_913_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/ptr_deref_913_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/ptr_deref_913_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/ptr_deref_913_Split/split_ack
      -- CP-element group 123: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/word_0/rr
      -- 
    rr_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(123), ack => ptr_deref_913_store_0_req_0); -- 
    convolution3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(90) & convolution3D_CP_1129_elements(94) & convolution3D_CP_1129_elements(98) & convolution3D_CP_1129_elements(102) & convolution3D_CP_1129_elements(106) & convolution3D_CP_1129_elements(110) & convolution3D_CP_1129_elements(114) & convolution3D_CP_1129_elements(118) & convolution3D_CP_1129_elements(122);
      gj_convolution3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/word_0/ra
      -- 
    ra_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_913_store_0_ack_0, ack => convolution3D_CP_1129_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	275 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/word_0/ca
      -- 
    ca_2128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_913_store_0_ack_1, ack => convolution3D_CP_1129_elements(125)); -- 
    -- CP-element group 126:  branch  join  transition  place  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	87 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926__exit__
      -- CP-element group 126: 	 branch_block_stmt_454/if_stmt_927__entry__
      -- CP-element group 126: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/$exit
      -- CP-element group 126: 	 branch_block_stmt_454/if_stmt_927_dead_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_454/if_stmt_927_eval_test/$entry
      -- CP-element group 126: 	 branch_block_stmt_454/if_stmt_927_eval_test/$exit
      -- CP-element group 126: 	 branch_block_stmt_454/if_stmt_927_eval_test/branch_req
      -- CP-element group 126: 	 branch_block_stmt_454/R_exitcond33_928_place
      -- CP-element group 126: 	 branch_block_stmt_454/if_stmt_927_if_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_454/if_stmt_927_else_link/$entry
      -- 
    branch_req_2136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(126), ack => if_stmt_927_branch_req_0); -- 
    convolution3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(87) & convolution3D_CP_1129_elements(125);
      gj_convolution3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	277 
    -- CP-element group 127: 	278 
    -- CP-element group 127:  members (24) 
      -- CP-element group 127: 	 branch_block_stmt_454/merge_stmt_933__exit__
      -- CP-element group 127: 	 branch_block_stmt_454/assign_stmt_940_to_assign_stmt_955__entry__
      -- CP-element group 127: 	 branch_block_stmt_454/assign_stmt_940_to_assign_stmt_955__exit__
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 127: 	 branch_block_stmt_454/if_stmt_927_if_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_454/if_stmt_927_if_link/if_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 127: 	 branch_block_stmt_454/assign_stmt_940_to_assign_stmt_955/$entry
      -- CP-element group 127: 	 branch_block_stmt_454/assign_stmt_940_to_assign_stmt_955/$exit
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/$entry
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_454/merge_stmt_933_PhiReqMerge
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/$entry
      -- CP-element group 127: 	 branch_block_stmt_454/merge_stmt_933_PhiAck/dummy
      -- CP-element group 127: 	 branch_block_stmt_454/merge_stmt_933_PhiAck/$exit
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/SplitProtocol/Update/cr
      -- CP-element group 127: 	 branch_block_stmt_454/merge_stmt_933_PhiAck/$entry
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/SplitProtocol/Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/SplitProtocol/Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/SplitProtocol/Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/SplitProtocol/$entry
      -- 
    if_choice_transition_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_927_branch_ack_1, ack => convolution3D_CP_1129_elements(127)); -- 
    cr_3409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(127), ack => type_cast_961_inst_req_1); -- 
    rr_3404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(127), ack => type_cast_961_inst_req_0); -- 
    -- CP-element group 128:  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	271 
    -- CP-element group 128: 	272 
    -- CP-element group 128:  members (12) 
      -- CP-element group 128: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/$entry
      -- CP-element group 128: 	 branch_block_stmt_454/if_stmt_927_else_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_454/if_stmt_927_else_link/else_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_454/forx_xbody_forx_xbody
      -- CP-element group 128: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/SplitProtocol/Update/cr
      -- CP-element group 128: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/$entry
      -- CP-element group 128: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_927_branch_ack_0, ack => convolution3D_CP_1129_elements(128)); -- 
    cr_3355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(128), ack => type_cast_767_inst_req_1); -- 
    rr_3350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(128), ack => type_cast_767_inst_req_0); -- 
    -- CP-element group 129:  transition  place  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	281 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	300 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_454/if_stmt_978_if_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_454/if_stmt_978_if_link/if_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_454/forx_xend_ifx_xend
      -- CP-element group 129: 	 branch_block_stmt_454/forx_xend_ifx_xend_PhiReq/$exit
      -- CP-element group 129: 	 branch_block_stmt_454/forx_xend_ifx_xend_PhiReq/$entry
      -- 
    if_choice_transition_2166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_978_branch_ack_1, ack => convolution3D_CP_1129_elements(129)); -- 
    -- CP-element group 130:  merge  fork  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	281 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	282 
    -- CP-element group 130: 	283 
    -- CP-element group 130:  members (20) 
      -- CP-element group 130: 	 branch_block_stmt_454/merge_stmt_984__exit__
      -- CP-element group 130: 	 branch_block_stmt_454/assign_stmt_990_to_assign_stmt_996__entry__
      -- CP-element group 130: 	 branch_block_stmt_454/assign_stmt_990_to_assign_stmt_996__exit__
      -- CP-element group 130: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 130: 	 branch_block_stmt_454/if_stmt_978_else_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_454/if_stmt_978_else_link/else_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_454/forx_xend_bbx_xnphx_xi
      -- CP-element group 130: 	 branch_block_stmt_454/assign_stmt_990_to_assign_stmt_996/$entry
      -- CP-element group 130: 	 branch_block_stmt_454/assign_stmt_990_to_assign_stmt_996/$exit
      -- CP-element group 130: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/$entry
      -- CP-element group 130: 	 branch_block_stmt_454/merge_stmt_984_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/$entry
      -- CP-element group 130: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_454/merge_stmt_984_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_454/merge_stmt_984_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_454/merge_stmt_984_PhiAck/$entry
      -- CP-element group 130: 	 branch_block_stmt_454/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_454/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- 
    else_choice_transition_2170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_978_branch_ack_0, ack => convolution3D_CP_1129_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	295 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_update_start_
      -- CP-element group 131: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_Update/cr
      -- 
    ra_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1027_inst_ack_0, ack => convolution3D_CP_1129_elements(131)); -- 
    cr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(131), ack => RPIPE_maxpool_input_pipe_1027_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_Sample/rr
      -- 
    ca_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1027_inst_ack_1, ack => convolution3D_CP_1129_elements(132)); -- 
    rr_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(132), ack => type_cast_1031_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_Sample/ra
      -- 
    ra_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1031_inst_ack_0, ack => convolution3D_CP_1129_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	295 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_Update/ca
      -- 
    ca_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1031_inst_ack_1, ack => convolution3D_CP_1129_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	295 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_sample_completed_
      -- 
    ra_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1046_inst_ack_0, ack => convolution3D_CP_1129_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	295 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_Update/$exit
      -- 
    ca_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1046_inst_ack_1, ack => convolution3D_CP_1129_elements(136)); -- 
    -- CP-element group 137:  branch  join  transition  place  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (10) 
      -- CP-element group 137: 	 branch_block_stmt_454/if_stmt_1053_else_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052__exit__
      -- CP-element group 137: 	 branch_block_stmt_454/if_stmt_1053__entry__
      -- CP-element group 137: 	 branch_block_stmt_454/if_stmt_1053_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_454/if_stmt_1053_eval_test/branch_req
      -- CP-element group 137: 	 branch_block_stmt_454/R_cmpx_xi_1054_place
      -- CP-element group 137: 	 branch_block_stmt_454/if_stmt_1053_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_454/if_stmt_1053_eval_test/$entry
      -- CP-element group 137: 	 branch_block_stmt_454/if_stmt_1053_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/$exit
      -- 
    branch_req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(137), ack => if_stmt_1053_branch_req_0); -- 
    convolution3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(134) & convolution3D_CP_1129_elements(136);
      gj_convolution3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	285 
    -- CP-element group 138: 	286 
    -- CP-element group 138: 	288 
    -- CP-element group 138: 	289 
    -- CP-element group 138:  members (20) 
      -- CP-element group 138: 	 branch_block_stmt_454/if_stmt_1053_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/if_stmt_1053_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/$entry
      -- 
    if_choice_transition_2233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1053_branch_ack_1, ack => convolution3D_CP_1129_elements(138)); -- 
    rr_3466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(138), ack => type_cast_1005_inst_req_0); -- 
    cr_3471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(138), ack => type_cast_1005_inst_req_1); -- 
    cr_3494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(138), ack => type_cast_1012_inst_req_1); -- 
    rr_3489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(138), ack => type_cast_1012_inst_req_0); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	296 
    -- CP-element group 139: 	297 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_454/if_stmt_1053_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_454/if_stmt_1053_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 139: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/SplitProtocol/Update/cr
      -- CP-element group 139: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/$entry
      -- CP-element group 139: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/$entry
      -- CP-element group 139: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- 
    else_choice_transition_2237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1053_branch_ack_0, ack => convolution3D_CP_1129_elements(139)); -- 
    cr_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(139), ack => type_cast_1063_inst_req_1); -- 
    rr_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(139), ack => type_cast_1063_inst_req_0); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	299 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	146 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_final_index_sum_regn_sample_complete
      -- CP-element group 140: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_final_index_sum_regn_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_final_index_sum_regn_Sample/ack
      -- 
    ack_2268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1092_index_offset_ack_0, ack => convolution3D_CP_1129_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	299 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (11) 
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_final_index_sum_regn_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_request/$entry
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_request/req
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_offset_calculated
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_final_index_sum_regn_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_root_address_calculated
      -- 
    ack_2273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1092_index_offset_ack_1, ack => convolution3D_CP_1129_elements(141)); -- 
    req_2282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(141), ack => addr_of_1093_final_reg_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_request/$exit
      -- CP-element group 142: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_request/ack
      -- 
    ack_2283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1093_final_reg_ack_0, ack => convolution3D_CP_1129_elements(142)); -- 
    -- CP-element group 143:  join  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	299 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (28) 
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/word_access_start/word_0/rr
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/ptr_deref_1096_Split/split_ack
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/ptr_deref_1096_Split/split_req
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/ptr_deref_1096_Split/$exit
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/ptr_deref_1096_Split/$entry
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_word_addrgen/root_register_ack
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_word_addrgen/root_register_req
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_word_addrgen/$exit
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_word_addrgen/$entry
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_base_addr_resize/base_resize_ack
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_base_addr_resize/base_resize_req
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_base_addr_resize/$exit
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_base_addr_resize/$entry
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_base_address_resized
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_word_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_base_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_complete/ack
      -- CP-element group 143: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_complete/$exit
      -- 
    ack_2288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1093_final_reg_ack_1, ack => convolution3D_CP_1129_elements(143)); -- 
    rr_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(143), ack => ptr_deref_1096_store_0_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/word_access_start/word_0/ra
      -- CP-element group 144: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_sample_completed_
      -- 
    ra_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1096_store_0_ack_0, ack => convolution3D_CP_1129_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	299 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Update/word_access_complete/word_0/ca
      -- CP-element group 145: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Update/word_access_complete/word_0/$exit
      -- 
    ca_2338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1096_store_0_ack_1, ack => convolution3D_CP_1129_elements(145)); -- 
    -- CP-element group 146:  join  transition  place  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	140 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	300 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098__exit__
      -- CP-element group 146: 	 branch_block_stmt_454/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 146: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/$exit
      -- CP-element group 146: 	 branch_block_stmt_454/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- CP-element group 146: 	 branch_block_stmt_454/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- 
    convolution3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(140) & convolution3D_CP_1129_elements(145);
      gj_convolution3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	300 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_sample_completed_
      -- 
    ra_2350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1103_inst_ack_0, ack => convolution3D_CP_1129_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	300 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	155 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_update_completed_
      -- 
    ca_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1103_inst_ack_1, ack => convolution3D_CP_1129_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	300 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_Sample/$exit
      -- 
    ra_2364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1107_inst_ack_0, ack => convolution3D_CP_1129_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	300 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	155 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_update_completed_
      -- 
    ca_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1107_inst_ack_1, ack => convolution3D_CP_1129_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	300 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_sample_completed_
      -- 
    ra_2378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_0, ack => convolution3D_CP_1129_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	300 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	155 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_update_completed_
      -- 
    ca_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_1, ack => convolution3D_CP_1129_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	300 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_sample_completed_
      -- 
    ra_2392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1115_inst_ack_0, ack => convolution3D_CP_1129_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	300 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_update_completed_
      -- 
    ca_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1115_inst_ack_1, ack => convolution3D_CP_1129_elements(154)); -- 
    -- CP-element group 155:  branch  join  transition  place  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	148 
    -- CP-element group 155: 	150 
    -- CP-element group 155: 	152 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (10) 
      -- CP-element group 155: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152__exit__
      -- CP-element group 155: 	 branch_block_stmt_454/if_stmt_1153__entry__
      -- CP-element group 155: 	 branch_block_stmt_454/R_cmp161321_1154_place
      -- CP-element group 155: 	 branch_block_stmt_454/if_stmt_1153_else_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_454/if_stmt_1153_if_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_454/if_stmt_1153_eval_test/branch_req
      -- CP-element group 155: 	 branch_block_stmt_454/if_stmt_1153_eval_test/$exit
      -- CP-element group 155: 	 branch_block_stmt_454/if_stmt_1153_eval_test/$entry
      -- CP-element group 155: 	 branch_block_stmt_454/if_stmt_1153_dead_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/$exit
      -- 
    branch_req_2405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(155), ack => if_stmt_1153_branch_req_0); -- 
    convolution3D_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(148) & convolution3D_CP_1129_elements(150) & convolution3D_CP_1129_elements(152) & convolution3D_CP_1129_elements(154);
      gj_convolution3D_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: 	159 
    -- CP-element group 156: 	160 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	162 
    -- CP-element group 156: 	163 
    -- CP-element group 156: 	164 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	168 
    -- CP-element group 156: 	170 
    -- CP-element group 156:  members (42) 
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/merge_stmt_1159_PhiReqMerge
      -- CP-element group 156: 	 branch_block_stmt_454/ifx_xend_bbx_xnph
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_update_start_
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_454/merge_stmt_1159__exit__
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230__entry__
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_update_start_
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/merge_stmt_1159_PhiAck/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_454/if_stmt_1153_if_link/if_choice_transition
      -- CP-element group 156: 	 branch_block_stmt_454/if_stmt_1153_if_link/$exit
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_update_start_
      -- CP-element group 156: 	 branch_block_stmt_454/merge_stmt_1159_PhiAck/$exit
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_update_start_
      -- CP-element group 156: 	 branch_block_stmt_454/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_454/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_update_start_
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_update_start_
      -- CP-element group 156: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_454/merge_stmt_1159_PhiAck/dummy
      -- 
    if_choice_transition_2410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1153_branch_ack_1, ack => convolution3D_CP_1129_elements(156)); -- 
    rr_2427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1174_inst_req_0); -- 
    cr_2432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1174_inst_req_1); -- 
    cr_2474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1196_inst_req_1); -- 
    rr_2469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1196_inst_req_0); -- 
    cr_2460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1187_inst_req_1); -- 
    rr_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1187_inst_req_0); -- 
    cr_2502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1210_inst_req_1); -- 
    cr_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1178_inst_req_1); -- 
    rr_2441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1178_inst_req_0); -- 
    cr_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1205_inst_req_1); -- 
    -- CP-element group 157:  transition  place  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	310 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_454/ifx_xend_forx_xend215
      -- CP-element group 157: 	 branch_block_stmt_454/if_stmt_1153_else_link/else_choice_transition
      -- CP-element group 157: 	 branch_block_stmt_454/if_stmt_1153_else_link/$exit
      -- CP-element group 157: 	 branch_block_stmt_454/ifx_xend_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$entry
      -- CP-element group 157: 	 branch_block_stmt_454/ifx_xend_forx_xend215_PhiReq/phi_stmt_1427/$entry
      -- CP-element group 157: 	 branch_block_stmt_454/ifx_xend_forx_xend215_PhiReq/$entry
      -- 
    else_choice_transition_2414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1153_branch_ack_0, ack => convolution3D_CP_1129_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_sample_completed_
      -- 
    ra_2428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_0, ack => convolution3D_CP_1129_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	156 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	166 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1174_Update/ca
      -- 
    ca_2433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_1, ack => convolution3D_CP_1129_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	156 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_Sample/ra
      -- CP-element group 160: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_sample_completed_
      -- 
    ra_2442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1178_inst_ack_0, ack => convolution3D_CP_1129_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	166 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_Update/ca
      -- CP-element group 161: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1178_update_completed_
      -- 
    ca_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1178_inst_ack_1, ack => convolution3D_CP_1129_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	156 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_Sample/ra
      -- CP-element group 162: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_sample_completed_
      -- 
    ra_2456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1187_inst_ack_0, ack => convolution3D_CP_1129_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	156 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	166 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_Update/ca
      -- CP-element group 163: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1187_update_completed_
      -- 
    ca_2461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1187_inst_ack_1, ack => convolution3D_CP_1129_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	156 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_Sample/ra
      -- CP-element group 164: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_sample_completed_
      -- 
    ra_2470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1196_inst_ack_0, ack => convolution3D_CP_1129_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	156 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_Update/ca
      -- CP-element group 165: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1196_update_completed_
      -- 
    ca_2475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1196_inst_ack_1, ack => convolution3D_CP_1129_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	159 
    -- CP-element group 166: 	161 
    -- CP-element group 166: 	163 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_sample_start_
      -- 
    rr_2483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(166), ack => type_cast_1205_inst_req_0); -- 
    convolution3D_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(159) & convolution3D_CP_1129_elements(161) & convolution3D_CP_1129_elements(163) & convolution3D_CP_1129_elements(165);
      gj_convolution3D_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_sample_completed_
      -- 
    ra_2484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1205_inst_ack_0, ack => convolution3D_CP_1129_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	156 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_Sample/rr
      -- CP-element group 168: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1205_Update/ca
      -- 
    ca_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1205_inst_ack_1, ack => convolution3D_CP_1129_elements(168)); -- 
    rr_2497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(168), ack => type_cast_1210_inst_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_Sample/ra
      -- CP-element group 169: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_sample_completed_
      -- 
    ra_2498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1210_inst_ack_0, ack => convolution3D_CP_1129_elements(169)); -- 
    -- CP-element group 170:  transition  place  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	156 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	301 
    -- CP-element group 170:  members (9) 
      -- CP-element group 170: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230__exit__
      -- CP-element group 170: 	 branch_block_stmt_454/bbx_xnph_forx_xbody163
      -- CP-element group 170: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/$exit
      -- CP-element group 170: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_Update/ca
      -- CP-element group 170: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_454/assign_stmt_1165_to_assign_stmt_1230/type_cast_1210_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_454/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/$entry
      -- CP-element group 170: 	 branch_block_stmt_454/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1233/$entry
      -- CP-element group 170: 	 branch_block_stmt_454/bbx_xnph_forx_xbody163_PhiReq/$entry
      -- 
    ca_2503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1210_inst_ack_1, ack => convolution3D_CP_1129_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	306 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	210 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_final_index_sum_regn_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_final_index_sum_regn_sample_complete
      -- CP-element group 171: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_final_index_sum_regn_Sample/ack
      -- 
    ack_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1245_index_offset_ack_0, ack => convolution3D_CP_1129_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	306 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (11) 
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_final_index_sum_regn_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_request/$entry
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_request/req
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_final_index_sum_regn_Update/ack
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_offset_calculated
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_sample_start_
      -- 
    ack_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1245_index_offset_ack_1, ack => convolution3D_CP_1129_elements(172)); -- 
    req_2546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(172), ack => addr_of_1246_final_reg_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_request/$exit
      -- CP-element group 173: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_request/ack
      -- 
    ack_2547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1246_final_reg_ack_0, ack => convolution3D_CP_1129_elements(173)); -- 
    -- CP-element group 174:  fork  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	306 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	207 
    -- CP-element group 174:  members (19) 
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_complete/$exit
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_complete/ack
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_base_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_word_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_root_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_base_address_resized
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_base_addr_resize/$entry
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_base_addr_resize/$exit
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_base_addr_resize/base_resize_req
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_base_addr_resize/base_resize_ack
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_base_plus_offset/$entry
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_base_plus_offset/$exit
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_base_plus_offset/sum_rename_req
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_base_plus_offset/sum_rename_ack
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_word_addrgen/$entry
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_word_addrgen/$exit
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_word_addrgen/root_register_req
      -- CP-element group 174: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_word_addrgen/root_register_ack
      -- 
    ack_2552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1246_final_reg_ack_1, ack => convolution3D_CP_1129_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	306 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_update_start_
      -- CP-element group 175: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_sample_completed_
      -- 
    ra_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1249_inst_ack_0, ack => convolution3D_CP_1129_elements(175)); -- 
    cr_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(175), ack => RPIPE_maxpool_input_pipe_1249_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_Sample/rr
      -- 
    ca_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1249_inst_ack_1, ack => convolution3D_CP_1129_elements(176)); -- 
    rr_2574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(176), ack => type_cast_1253_inst_req_0); -- 
    rr_2588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(176), ack => RPIPE_maxpool_input_pipe_1262_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_sample_completed_
      -- 
    ra_2575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1253_inst_ack_0, ack => convolution3D_CP_1129_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	306 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	207 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_update_completed_
      -- 
    ca_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1253_inst_ack_1, ack => convolution3D_CP_1129_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_update_start_
      -- CP-element group 179: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_Update/cr
      -- CP-element group 179: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_Sample/ra
      -- 
    ra_2589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1262_inst_ack_0, ack => convolution3D_CP_1129_elements(179)); -- 
    cr_2593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(179), ack => RPIPE_maxpool_input_pipe_1262_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1262_Update/$exit
      -- 
    ca_2594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1262_inst_ack_1, ack => convolution3D_CP_1129_elements(180)); -- 
    rr_2602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(180), ack => type_cast_1266_inst_req_0); -- 
    rr_2616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(180), ack => RPIPE_maxpool_input_pipe_1280_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_sample_completed_
      -- 
    ra_2603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_0, ack => convolution3D_CP_1129_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	306 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	207 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_update_completed_
      -- 
    ca_2608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_1, ack => convolution3D_CP_1129_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_Update/cr
      -- CP-element group 183: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_update_start_
      -- CP-element group 183: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_sample_completed_
      -- 
    ra_2617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1280_inst_ack_0, ack => convolution3D_CP_1129_elements(183)); -- 
    cr_2621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(183), ack => RPIPE_maxpool_input_pipe_1280_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1280_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_Sample/rr
      -- 
    ca_2622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1280_inst_ack_1, ack => convolution3D_CP_1129_elements(184)); -- 
    rr_2630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(184), ack => type_cast_1284_inst_req_0); -- 
    rr_2644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(184), ack => RPIPE_maxpool_input_pipe_1298_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_Sample/$exit
      -- 
    ra_2631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_0, ack => convolution3D_CP_1129_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	306 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	207 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_Update/$exit
      -- 
    ca_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_1, ack => convolution3D_CP_1129_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_Update/cr
      -- CP-element group 187: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_update_start_
      -- CP-element group 187: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_sample_completed_
      -- 
    ra_2645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1298_inst_ack_0, ack => convolution3D_CP_1129_elements(187)); -- 
    cr_2649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(187), ack => RPIPE_maxpool_input_pipe_1298_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1298_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_Sample/$entry
      -- 
    ca_2650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1298_inst_ack_1, ack => convolution3D_CP_1129_elements(188)); -- 
    rr_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(188), ack => type_cast_1302_inst_req_0); -- 
    rr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(188), ack => RPIPE_maxpool_input_pipe_1316_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_sample_completed_
      -- 
    ra_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1302_inst_ack_0, ack => convolution3D_CP_1129_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	306 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	207 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_Update/ca
      -- 
    ca_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1302_inst_ack_1, ack => convolution3D_CP_1129_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_update_start_
      -- CP-element group 191: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_Update/cr
      -- CP-element group 191: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_Sample/$exit
      -- 
    ra_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1316_inst_ack_0, ack => convolution3D_CP_1129_elements(191)); -- 
    cr_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(191), ack => RPIPE_maxpool_input_pipe_1316_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1316_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_sample_start_
      -- 
    ca_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1316_inst_ack_1, ack => convolution3D_CP_1129_elements(192)); -- 
    rr_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(192), ack => type_cast_1320_inst_req_0); -- 
    rr_2700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(192), ack => RPIPE_maxpool_input_pipe_1334_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_Sample/$exit
      -- 
    ra_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_0, ack => convolution3D_CP_1129_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	306 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	207 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_Update/$exit
      -- 
    ca_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_1, ack => convolution3D_CP_1129_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_update_start_
      -- CP-element group 195: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_Update/cr
      -- 
    ra_2701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1334_inst_ack_0, ack => convolution3D_CP_1129_elements(195)); -- 
    cr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(195), ack => RPIPE_maxpool_input_pipe_1334_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1334_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_Sample/rr
      -- 
    ca_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1334_inst_ack_1, ack => convolution3D_CP_1129_elements(196)); -- 
    rr_2714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(196), ack => type_cast_1338_inst_req_0); -- 
    rr_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(196), ack => RPIPE_maxpool_input_pipe_1352_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_Sample/ra
      -- 
    ra_2715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_0, ack => convolution3D_CP_1129_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	306 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	207 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_Update/ca
      -- 
    ca_2720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_1, ack => convolution3D_CP_1129_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_update_start_
      -- CP-element group 199: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_Update/cr
      -- 
    ra_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1352_inst_ack_0, ack => convolution3D_CP_1129_elements(199)); -- 
    cr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(199), ack => RPIPE_maxpool_input_pipe_1352_inst_req_1); -- 
    -- CP-element group 200:  fork  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200: 	203 
    -- CP-element group 200:  members (9) 
      -- CP-element group 200: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1352_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_Sample/rr
      -- 
    ca_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1352_inst_ack_1, ack => convolution3D_CP_1129_elements(200)); -- 
    rr_2742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(200), ack => type_cast_1356_inst_req_0); -- 
    rr_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(200), ack => RPIPE_maxpool_input_pipe_1370_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_Sample/ra
      -- 
    ra_2743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_0, ack => convolution3D_CP_1129_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	306 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	207 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_Update/ca
      -- 
    ca_2748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_1, ack => convolution3D_CP_1129_elements(202)); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	200 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_update_start_
      -- CP-element group 203: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_Sample/ra
      -- CP-element group 203: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_Update/cr
      -- 
    ra_2757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1370_inst_ack_0, ack => convolution3D_CP_1129_elements(203)); -- 
    cr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(203), ack => RPIPE_maxpool_input_pipe_1370_inst_req_1); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1370_Update/ca
      -- CP-element group 204: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_Sample/rr
      -- 
    ca_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1370_inst_ack_1, ack => convolution3D_CP_1129_elements(204)); -- 
    rr_2770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(204), ack => type_cast_1374_inst_req_0); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_Sample/ra
      -- 
    ra_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1374_inst_ack_0, ack => convolution3D_CP_1129_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	306 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_Update/ca
      -- 
    ca_2776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1374_inst_ack_1, ack => convolution3D_CP_1129_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	174 
    -- CP-element group 207: 	178 
    -- CP-element group 207: 	182 
    -- CP-element group 207: 	186 
    -- CP-element group 207: 	190 
    -- CP-element group 207: 	194 
    -- CP-element group 207: 	198 
    -- CP-element group 207: 	202 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/ptr_deref_1382_Split/$entry
      -- CP-element group 207: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/ptr_deref_1382_Split/$exit
      -- CP-element group 207: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/ptr_deref_1382_Split/split_req
      -- CP-element group 207: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/ptr_deref_1382_Split/split_ack
      -- CP-element group 207: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/word_access_start/$entry
      -- CP-element group 207: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/word_access_start/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/word_access_start/word_0/rr
      -- 
    rr_2814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(207), ack => ptr_deref_1382_store_0_req_0); -- 
    convolution3D_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(174) & convolution3D_CP_1129_elements(178) & convolution3D_CP_1129_elements(182) & convolution3D_CP_1129_elements(186) & convolution3D_CP_1129_elements(190) & convolution3D_CP_1129_elements(194) & convolution3D_CP_1129_elements(198) & convolution3D_CP_1129_elements(202) & convolution3D_CP_1129_elements(206);
      gj_convolution3D_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/word_access_start/$exit
      -- CP-element group 208: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/word_access_start/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Sample/word_access_start/word_0/ra
      -- 
    ra_2815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_store_0_ack_0, ack => convolution3D_CP_1129_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	306 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Update/word_access_complete/$exit
      -- CP-element group 209: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Update/word_access_complete/word_0/$exit
      -- CP-element group 209: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Update/word_access_complete/word_0/ca
      -- 
    ca_2826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_store_0_ack_1, ack => convolution3D_CP_1129_elements(209)); -- 
    -- CP-element group 210:  branch  join  transition  place  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	171 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (10) 
      -- CP-element group 210: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395__exit__
      -- CP-element group 210: 	 branch_block_stmt_454/if_stmt_1396__entry__
      -- CP-element group 210: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/$exit
      -- CP-element group 210: 	 branch_block_stmt_454/if_stmt_1396_dead_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_454/if_stmt_1396_eval_test/$entry
      -- CP-element group 210: 	 branch_block_stmt_454/if_stmt_1396_eval_test/$exit
      -- CP-element group 210: 	 branch_block_stmt_454/if_stmt_1396_eval_test/branch_req
      -- CP-element group 210: 	 branch_block_stmt_454/R_exitcond_1397_place
      -- CP-element group 210: 	 branch_block_stmt_454/if_stmt_1396_if_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_454/if_stmt_1396_else_link/$entry
      -- 
    branch_req_2834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(210), ack => if_stmt_1396_branch_req_0); -- 
    convolution3D_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(171) & convolution3D_CP_1129_elements(209);
      gj_convolution3D_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	307 
    -- CP-element group 211: 	308 
    -- CP-element group 211:  members (24) 
      -- CP-element group 211: 	 branch_block_stmt_454/merge_stmt_1402_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_454/merge_stmt_1402_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_454/merge_stmt_1402_PhiReqMerge
      -- CP-element group 211: 	 branch_block_stmt_454/merge_stmt_1402__exit__
      -- CP-element group 211: 	 branch_block_stmt_454/assign_stmt_1409_to_assign_stmt_1424__entry__
      -- CP-element group 211: 	 branch_block_stmt_454/assign_stmt_1409_to_assign_stmt_1424__exit__
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215
      -- CP-element group 211: 	 branch_block_stmt_454/merge_stmt_1402_PhiAck/dummy
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_454/if_stmt_1396_if_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_454/if_stmt_1396_if_link/if_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge
      -- CP-element group 211: 	 branch_block_stmt_454/assign_stmt_1409_to_assign_stmt_1424/$entry
      -- CP-element group 211: 	 branch_block_stmt_454/assign_stmt_1409_to_assign_stmt_1424/$exit
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$entry
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Update/cr
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/$entry
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/$entry
      -- CP-element group 211: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/$entry
      -- 
    if_choice_transition_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1396_branch_ack_1, ack => convolution3D_CP_1129_elements(211)); -- 
    cr_3638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(211), ack => type_cast_1430_inst_req_1); -- 
    rr_3633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(211), ack => type_cast_1430_inst_req_0); -- 
    -- CP-element group 212:  fork  transition  place  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	302 
    -- CP-element group 212: 	303 
    -- CP-element group 212:  members (12) 
      -- CP-element group 212: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/SplitProtocol/Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/SplitProtocol/Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/SplitProtocol/Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/SplitProtocol/$entry
      -- CP-element group 212: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/$entry
      -- CP-element group 212: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/$entry
      -- CP-element group 212: 	 branch_block_stmt_454/if_stmt_1396_else_link/$exit
      -- CP-element group 212: 	 branch_block_stmt_454/if_stmt_1396_else_link/else_choice_transition
      -- CP-element group 212: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163
      -- CP-element group 212: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1396_branch_ack_0, ack => convolution3D_CP_1129_elements(212)); -- 
    rr_3590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(212), ack => type_cast_1239_inst_req_0); -- 
    cr_3595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(212), ack => type_cast_1239_inst_req_1); -- 
    -- CP-element group 213:  transition  place  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	312 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	331 
    -- CP-element group 213:  members (5) 
      -- CP-element group 213: 	 branch_block_stmt_454/if_stmt_1447_if_link/$exit
      -- CP-element group 213: 	 branch_block_stmt_454/if_stmt_1447_if_link/if_choice_transition
      -- CP-element group 213: 	 branch_block_stmt_454/forx_xend215_ifx_xend227
      -- CP-element group 213: 	 branch_block_stmt_454/forx_xend215_ifx_xend227_PhiReq/$entry
      -- CP-element group 213: 	 branch_block_stmt_454/forx_xend215_ifx_xend227_PhiReq/$exit
      -- 
    if_choice_transition_2864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1447_branch_ack_1, ack => convolution3D_CP_1129_elements(213)); -- 
    -- CP-element group 214:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	312 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (18) 
      -- CP-element group 214: 	 branch_block_stmt_454/merge_stmt_1453_PhiReqMerge
      -- CP-element group 214: 	 branch_block_stmt_454/merge_stmt_1453__exit__
      -- CP-element group 214: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469__entry__
      -- CP-element group 214: 	 branch_block_stmt_454/forx_xend215_bbx_xnphx_xi298_PhiReq/$exit
      -- CP-element group 214: 	 branch_block_stmt_454/if_stmt_1447_else_link/$exit
      -- CP-element group 214: 	 branch_block_stmt_454/if_stmt_1447_else_link/else_choice_transition
      -- CP-element group 214: 	 branch_block_stmt_454/forx_xend215_bbx_xnphx_xi298
      -- CP-element group 214: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/$entry
      -- CP-element group 214: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_update_start_
      -- CP-element group 214: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_Sample/rr
      -- CP-element group 214: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_Update/cr
      -- CP-element group 214: 	 branch_block_stmt_454/merge_stmt_1453_PhiAck/dummy
      -- CP-element group 214: 	 branch_block_stmt_454/merge_stmt_1453_PhiAck/$exit
      -- CP-element group 214: 	 branch_block_stmt_454/merge_stmt_1453_PhiAck/$entry
      -- CP-element group 214: 	 branch_block_stmt_454/forx_xend215_bbx_xnphx_xi298_PhiReq/$entry
      -- 
    else_choice_transition_2868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1447_branch_ack_0, ack => convolution3D_CP_1129_elements(214)); -- 
    rr_2881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(214), ack => type_cast_1462_inst_req_0); -- 
    cr_2886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(214), ack => type_cast_1462_inst_req_1); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_Sample/ra
      -- 
    ra_2882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1462_inst_ack_0, ack => convolution3D_CP_1129_elements(215)); -- 
    -- CP-element group 216:  fork  transition  place  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	313 
    -- CP-element group 216: 	314 
    -- CP-element group 216:  members (11) 
      -- CP-element group 216: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469__exit__
      -- CP-element group 216: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307
      -- CP-element group 216: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/$entry
      -- CP-element group 216: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/$entry
      -- CP-element group 216: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/$exit
      -- CP-element group 216: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_454/assign_stmt_1459_to_assign_stmt_1469/type_cast_1462_Update/ca
      -- CP-element group 216: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/$entry
      -- 
    ca_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1462_inst_ack_1, ack => convolution3D_CP_1129_elements(216)); -- 
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	326 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_update_start_
      -- CP-element group 217: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_Sample/ra
      -- CP-element group 217: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_Update/cr
      -- 
    ra_2899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1500_inst_ack_0, ack => convolution3D_CP_1129_elements(217)); -- 
    cr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(217), ack => RPIPE_maxpool_input_pipe_1500_inst_req_1); -- 
    -- CP-element group 218:  transition  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (6) 
      -- CP-element group 218: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_Update/ca
      -- CP-element group 218: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_Sample/rr
      -- 
    ca_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1500_inst_ack_1, ack => convolution3D_CP_1129_elements(218)); -- 
    rr_2912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(218), ack => type_cast_1504_inst_req_0); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_Sample/ra
      -- 
    ra_2913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1504_inst_ack_0, ack => convolution3D_CP_1129_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	326 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	223 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_Update/ca
      -- 
    ca_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1504_inst_ack_1, ack => convolution3D_CP_1129_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	326 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_Sample/ra
      -- 
    ra_2927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1519_inst_ack_0, ack => convolution3D_CP_1129_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	326 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_Update/ca
      -- 
    ca_2932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1519_inst_ack_1, ack => convolution3D_CP_1129_elements(222)); -- 
    -- CP-element group 223:  branch  join  transition  place  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	220 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (10) 
      -- CP-element group 223: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525__exit__
      -- CP-element group 223: 	 branch_block_stmt_454/if_stmt_1526__entry__
      -- CP-element group 223: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/$exit
      -- CP-element group 223: 	 branch_block_stmt_454/if_stmt_1526_dead_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_454/if_stmt_1526_eval_test/$entry
      -- CP-element group 223: 	 branch_block_stmt_454/if_stmt_1526_eval_test/$exit
      -- CP-element group 223: 	 branch_block_stmt_454/if_stmt_1526_eval_test/branch_req
      -- CP-element group 223: 	 branch_block_stmt_454/R_cmpx_xi306_1527_place
      -- CP-element group 223: 	 branch_block_stmt_454/if_stmt_1526_if_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_454/if_stmt_1526_else_link/$entry
      -- 
    branch_req_2940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(223), ack => if_stmt_1526_branch_req_0); -- 
    convolution3D_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(220) & convolution3D_CP_1129_elements(222);
      gj_convolution3D_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  place  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	316 
    -- CP-element group 224: 	317 
    -- CP-element group 224: 	319 
    -- CP-element group 224: 	320 
    -- CP-element group 224:  members (20) 
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/SplitProtocol/Update/cr
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_454/if_stmt_1526_if_link/$exit
      -- CP-element group 224: 	 branch_block_stmt_454/if_stmt_1526_if_link/if_choice_transition
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1526_branch_ack_1, ack => convolution3D_CP_1129_elements(224)); -- 
    cr_3711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(224), ack => type_cast_1478_inst_req_1); -- 
    rr_3706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(224), ack => type_cast_1478_inst_req_0); -- 
    rr_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(224), ack => type_cast_1485_inst_req_0); -- 
    cr_3734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(224), ack => type_cast_1485_inst_req_1); -- 
    -- CP-element group 225:  fork  transition  place  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	327 
    -- CP-element group 225: 	328 
    -- CP-element group 225:  members (12) 
      -- CP-element group 225: 	 branch_block_stmt_454/if_stmt_1526_else_link/$exit
      -- CP-element group 225: 	 branch_block_stmt_454/if_stmt_1526_else_link/else_choice_transition
      -- CP-element group 225: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315
      -- CP-element group 225: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/$entry
      -- CP-element group 225: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/$entry
      -- CP-element group 225: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/$entry
      -- CP-element group 225: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/$entry
      -- CP-element group 225: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/SplitProtocol/$entry
      -- CP-element group 225: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/SplitProtocol/Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/SplitProtocol/Sample/rr
      -- CP-element group 225: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/SplitProtocol/Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1526_branch_ack_0, ack => convolution3D_CP_1129_elements(225)); -- 
    rr_3765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(225), ack => type_cast_1536_inst_req_0); -- 
    cr_3770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(225), ack => type_cast_1536_inst_req_1); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	330 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	232 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_final_index_sum_regn_sample_complete
      -- CP-element group 226: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_final_index_sum_regn_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_final_index_sum_regn_Sample/ack
      -- 
    ack_2980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1565_index_offset_ack_0, ack => convolution3D_CP_1129_elements(226)); -- 
    -- CP-element group 227:  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	330 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (11) 
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_root_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_offset_calculated
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_final_index_sum_regn_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_final_index_sum_regn_Update/ack
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_base_plus_offset/$entry
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_base_plus_offset/$exit
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_base_plus_offset/sum_rename_req
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_base_plus_offset/sum_rename_ack
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_request/$entry
      -- CP-element group 227: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_request/req
      -- 
    ack_2985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1565_index_offset_ack_1, ack => convolution3D_CP_1129_elements(227)); -- 
    req_2994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(227), ack => addr_of_1566_final_reg_req_0); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_request/$exit
      -- CP-element group 228: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_request/ack
      -- 
    ack_2995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1566_final_reg_ack_0, ack => convolution3D_CP_1129_elements(228)); -- 
    -- CP-element group 229:  join  fork  transition  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	330 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (28) 
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_complete/$exit
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_complete/ack
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_base_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_word_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_root_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_base_address_resized
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_base_addr_resize/$entry
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_base_addr_resize/$exit
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_base_addr_resize/base_resize_req
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_base_addr_resize/base_resize_ack
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_base_plus_offset/$entry
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_base_plus_offset/$exit
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_base_plus_offset/sum_rename_req
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_base_plus_offset/sum_rename_ack
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_word_addrgen/$entry
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_word_addrgen/$exit
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_word_addrgen/root_register_req
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_word_addrgen/root_register_ack
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/ptr_deref_1569_Split/$entry
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/ptr_deref_1569_Split/$exit
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/ptr_deref_1569_Split/split_req
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/ptr_deref_1569_Split/split_ack
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/word_access_start/$entry
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/word_access_start/word_0/$entry
      -- CP-element group 229: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/word_access_start/word_0/rr
      -- 
    ack_3000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1566_final_reg_ack_1, ack => convolution3D_CP_1129_elements(229)); -- 
    rr_3038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(229), ack => ptr_deref_1569_store_0_req_0); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/word_access_start/$exit
      -- CP-element group 230: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/word_access_start/word_0/$exit
      -- CP-element group 230: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Sample/word_access_start/word_0/ra
      -- 
    ra_3039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1569_store_0_ack_0, ack => convolution3D_CP_1129_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	330 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (5) 
      -- CP-element group 231: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Update/word_access_complete/$exit
      -- CP-element group 231: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Update/word_access_complete/word_0/$exit
      -- CP-element group 231: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Update/word_access_complete/word_0/ca
      -- 
    ca_3050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1569_store_0_ack_1, ack => convolution3D_CP_1129_elements(231)); -- 
    -- CP-element group 232:  join  transition  place  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	226 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	331 
    -- CP-element group 232:  members (5) 
      -- CP-element group 232: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571__exit__
      -- CP-element group 232: 	 branch_block_stmt_454/getRemainingElementsx_xexit315_ifx_xend227
      -- CP-element group 232: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/$exit
      -- CP-element group 232: 	 branch_block_stmt_454/getRemainingElementsx_xexit315_ifx_xend227_PhiReq/$entry
      -- CP-element group 232: 	 branch_block_stmt_454/getRemainingElementsx_xexit315_ifx_xend227_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(226) & convolution3D_CP_1129_elements(231);
      gj_convolution3D_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	331 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_Sample/cra
      -- 
    cra_3062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1576_call_ack_0, ack => convolution3D_CP_1129_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	331 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	239 
    -- CP-element group 234: 	240 
    -- CP-element group 234: 	241 
    -- CP-element group 234: 	242 
    -- CP-element group 234: 	243 
    -- CP-element group 234: 	244 
    -- CP-element group 234:  members (28) 
      -- CP-element group 234: 	 branch_block_stmt_454/call_stmt_1576__exit__
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641__entry__
      -- CP-element group 234: 	 branch_block_stmt_454/call_stmt_1576/$exit
      -- CP-element group 234: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_Update/cca
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/$entry
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_update_start_
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_update_start_
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_update_start_
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_Update/cr
      -- 
    cca_3067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1576_call_ack_1, ack => convolution3D_CP_1129_elements(234)); -- 
    req_3078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => WPIPE_maxpool_output_pipe_1583_inst_req_0); -- 
    rr_3106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1616_inst_req_0); -- 
    cr_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1616_inst_req_1); -- 
    rr_3120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1626_inst_req_0); -- 
    cr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1626_inst_req_1); -- 
    rr_3134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1635_inst_req_0); -- 
    cr_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1635_inst_req_1); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_update_start_
      -- CP-element group 235: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_Update/req
      -- 
    ack_3079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1583_inst_ack_0, ack => convolution3D_CP_1129_elements(235)); -- 
    req_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(235), ack => WPIPE_maxpool_output_pipe_1583_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1583_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_Sample/req
      -- 
    ack_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1583_inst_ack_1, ack => convolution3D_CP_1129_elements(236)); -- 
    req_3092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(236), ack => WPIPE_maxpool_output_pipe_1587_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_update_start_
      -- CP-element group 237: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_Update/req
      -- 
    ack_3093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1587_inst_ack_0, ack => convolution3D_CP_1129_elements(237)); -- 
    req_3097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(237), ack => WPIPE_maxpool_output_pipe_1587_inst_req_1); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	245 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/WPIPE_maxpool_output_pipe_1587_Update/ack
      -- 
    ack_3098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1587_inst_ack_1, ack => convolution3D_CP_1129_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	234 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_Sample/ra
      -- 
    ra_3107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1616_inst_ack_0, ack => convolution3D_CP_1129_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	234 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	245 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1616_Update/ca
      -- 
    ca_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1616_inst_ack_1, ack => convolution3D_CP_1129_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	234 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_Sample/ra
      -- 
    ra_3121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1626_inst_ack_0, ack => convolution3D_CP_1129_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	234 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	245 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1626_Update/ca
      -- 
    ca_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1626_inst_ack_1, ack => convolution3D_CP_1129_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	234 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_Sample/ra
      -- 
    ra_3135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1635_inst_ack_0, ack => convolution3D_CP_1129_elements(243)); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	234 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/type_cast_1635_Update/ca
      -- 
    ca_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1635_inst_ack_1, ack => convolution3D_CP_1129_elements(244)); -- 
    -- CP-element group 245:  join  transition  place  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	238 
    -- CP-element group 245: 	240 
    -- CP-element group 245: 	242 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	332 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641__exit__
      -- CP-element group 245: 	 branch_block_stmt_454/ifx_xend227_whilex_xbody
      -- CP-element group 245: 	 branch_block_stmt_454/assign_stmt_1582_to_assign_stmt_1641/$exit
      -- CP-element group 245: 	 branch_block_stmt_454/ifx_xend227_whilex_xbody_PhiReq/$entry
      -- CP-element group 245: 	 branch_block_stmt_454/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1644/$entry
      -- CP-element group 245: 	 branch_block_stmt_454/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/$entry
      -- 
    convolution3D_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(238) & convolution3D_CP_1129_elements(240) & convolution3D_CP_1129_elements(242) & convolution3D_CP_1129_elements(244);
      gj_convolution3D_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	337 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_Sample/ra
      -- 
    ra_3152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1664_inst_ack_0, ack => convolution3D_CP_1129_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	337 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	254 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_Update/ca
      -- 
    ca_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1664_inst_ack_1, ack => convolution3D_CP_1129_elements(247)); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	337 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_update_start_
      -- CP-element group 248: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_Sample/ack
      -- CP-element group 248: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_Update/$entry
      -- CP-element group 248: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_Update/req
      -- 
    ack_3166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1666_inst_ack_0, ack => convolution3D_CP_1129_elements(248)); -- 
    req_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(248), ack => WPIPE_num_out_pipe_1666_inst_req_1); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	259 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_Update/ack
      -- 
    ack_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1666_inst_ack_1, ack => convolution3D_CP_1129_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	337 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_Sample/ra
      -- 
    ra_3180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1671_inst_ack_0, ack => convolution3D_CP_1129_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	337 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	254 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_Update/ca
      -- 
    ca_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1671_inst_ack_1, ack => convolution3D_CP_1129_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	337 
    -- CP-element group 252: successors 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_Sample/ra
      -- 
    ra_3194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1675_inst_ack_0, ack => convolution3D_CP_1129_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	337 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_Update/ca
      -- 
    ca_3199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1675_inst_ack_1, ack => convolution3D_CP_1129_elements(253)); -- 
    -- CP-element group 254:  join  transition  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	247 
    -- CP-element group 254: 	251 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_Sample/crr
      -- 
    crr_3207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(254), ack => call_stmt_1686_call_req_0); -- 
    convolution3D_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(247) & convolution3D_CP_1129_elements(251) & convolution3D_CP_1129_elements(253);
      gj_convolution3D_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_Sample/cra
      -- 
    cra_3208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1686_call_ack_0, ack => convolution3D_CP_1129_elements(255)); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	337 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	259 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_Update/cca
      -- 
    cca_3213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1686_call_ack_1, ack => convolution3D_CP_1129_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	337 
    -- CP-element group 257: successors 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_Sample/cra
      -- 
    cra_3222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1693_call_ack_0, ack => convolution3D_CP_1129_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	337 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_Update/cca
      -- 
    cca_3227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1693_call_ack_1, ack => convolution3D_CP_1129_elements(258)); -- 
    -- CP-element group 259:  branch  join  transition  place  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	249 
    -- CP-element group 259: 	256 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259: 	261 
    -- CP-element group 259:  members (10) 
      -- CP-element group 259: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704__exit__
      -- CP-element group 259: 	 branch_block_stmt_454/if_stmt_1705__entry__
      -- CP-element group 259: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/$exit
      -- CP-element group 259: 	 branch_block_stmt_454/if_stmt_1705_dead_link/$entry
      -- CP-element group 259: 	 branch_block_stmt_454/if_stmt_1705_eval_test/$entry
      -- CP-element group 259: 	 branch_block_stmt_454/if_stmt_1705_eval_test/$exit
      -- CP-element group 259: 	 branch_block_stmt_454/if_stmt_1705_eval_test/branch_req
      -- CP-element group 259: 	 branch_block_stmt_454/R_exitcond5_1706_place
      -- CP-element group 259: 	 branch_block_stmt_454/if_stmt_1705_if_link/$entry
      -- CP-element group 259: 	 branch_block_stmt_454/if_stmt_1705_else_link/$entry
      -- 
    branch_req_3235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(259), ack => if_stmt_1705_branch_req_0); -- 
    convolution3D_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(249) & convolution3D_CP_1129_elements(256) & convolution3D_CP_1129_elements(258);
      gj_convolution3D_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260: 	263 
    -- CP-element group 260:  members (18) 
      -- CP-element group 260: 	 branch_block_stmt_454/merge_stmt_1711__exit__
      -- CP-element group 260: 	 branch_block_stmt_454/assign_stmt_1716__entry__
      -- CP-element group 260: 	 branch_block_stmt_454/merge_stmt_1711_PhiReqMerge
      -- CP-element group 260: 	 branch_block_stmt_454/if_stmt_1705_if_link/$exit
      -- CP-element group 260: 	 branch_block_stmt_454/if_stmt_1705_if_link/if_choice_transition
      -- CP-element group 260: 	 branch_block_stmt_454/whilex_xbody_whilex_xend
      -- CP-element group 260: 	 branch_block_stmt_454/assign_stmt_1716/$entry
      -- CP-element group 260: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_update_start_
      -- CP-element group 260: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_Sample/rr
      -- CP-element group 260: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_Update/cr
      -- CP-element group 260: 	 branch_block_stmt_454/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 260: 	 branch_block_stmt_454/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 260: 	 branch_block_stmt_454/merge_stmt_1711_PhiAck/$entry
      -- CP-element group 260: 	 branch_block_stmt_454/merge_stmt_1711_PhiAck/$exit
      -- CP-element group 260: 	 branch_block_stmt_454/merge_stmt_1711_PhiAck/dummy
      -- 
    if_choice_transition_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1705_branch_ack_1, ack => convolution3D_CP_1129_elements(260)); -- 
    rr_3257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(260), ack => type_cast_1715_inst_req_0); -- 
    cr_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(260), ack => type_cast_1715_inst_req_1); -- 
    -- CP-element group 261:  fork  transition  place  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	259 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	333 
    -- CP-element group 261: 	334 
    -- CP-element group 261:  members (12) 
      -- CP-element group 261: 	 branch_block_stmt_454/if_stmt_1705_else_link/$exit
      -- CP-element group 261: 	 branch_block_stmt_454/if_stmt_1705_else_link/else_choice_transition
      -- CP-element group 261: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody
      -- CP-element group 261: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 261: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/$entry
      -- CP-element group 261: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/$entry
      -- CP-element group 261: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/$entry
      -- CP-element group 261: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/SplitProtocol/$entry
      -- CP-element group 261: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/SplitProtocol/Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/SplitProtocol/Sample/rr
      -- CP-element group 261: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/SplitProtocol/Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1705_branch_ack_0, ack => convolution3D_CP_1129_elements(261)); -- 
    rr_3818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(261), ack => type_cast_1647_inst_req_0); -- 
    cr_3823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(261), ack => type_cast_1647_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_sample_completed_
      -- CP-element group 262: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_Sample/ra
      -- 
    ra_3258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1715_inst_ack_0, ack => convolution3D_CP_1129_elements(262)); -- 
    -- CP-element group 263:  fork  transition  place  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	260 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263: 	265 
    -- CP-element group 263: 	267 
    -- CP-element group 263:  members (16) 
      -- CP-element group 263: 	 branch_block_stmt_454/assign_stmt_1716__exit__
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732__entry__
      -- CP-element group 263: 	 branch_block_stmt_454/assign_stmt_1716/$exit
      -- CP-element group 263: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_update_completed_
      -- CP-element group 263: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_454/assign_stmt_1716/type_cast_1715_Update/ca
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/$entry
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_update_start_
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_Sample/crr
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_Update/ccr
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_update_start_
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_Update/cr
      -- 
    ca_3263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1715_inst_ack_1, ack => convolution3D_CP_1129_elements(263)); -- 
    crr_3274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => call_stmt_1719_call_req_0); -- 
    ccr_3279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => call_stmt_1719_call_req_1); -- 
    cr_3293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => type_cast_1723_inst_req_1); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_Sample/cra
      -- 
    cra_3275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1719_call_ack_0, ack => convolution3D_CP_1129_elements(264)); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/call_stmt_1719_Update/cca
      -- CP-element group 265: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_Sample/rr
      -- 
    cca_3280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1719_call_ack_1, ack => convolution3D_CP_1129_elements(265)); -- 
    rr_3288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(265), ack => type_cast_1723_inst_req_0); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_Sample/ra
      -- 
    ra_3289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1723_inst_ack_0, ack => convolution3D_CP_1129_elements(266)); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	263 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/type_cast_1723_Update/ca
      -- CP-element group 267: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_Sample/req
      -- 
    ca_3294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1723_inst_ack_1, ack => convolution3D_CP_1129_elements(267)); -- 
    req_3302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(267), ack => WPIPE_elapsed_time_pipe_1730_inst_req_0); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_update_start_
      -- CP-element group 268: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_Sample/ack
      -- CP-element group 268: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_Update/$entry
      -- CP-element group 268: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_Update/req
      -- 
    ack_3303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1730_inst_ack_0, ack => convolution3D_CP_1129_elements(268)); -- 
    req_3307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(268), ack => WPIPE_elapsed_time_pipe_1730_inst_req_1); -- 
    -- CP-element group 269:  transition  place  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269:  members (16) 
      -- CP-element group 269: 	 $exit
      -- CP-element group 269: 	 branch_block_stmt_454/$exit
      -- CP-element group 269: 	 branch_block_stmt_454/branch_block_stmt_454__exit__
      -- CP-element group 269: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732__exit__
      -- CP-element group 269: 	 branch_block_stmt_454/return__
      -- CP-element group 269: 	 branch_block_stmt_454/merge_stmt_1735__exit__
      -- CP-element group 269: 	 branch_block_stmt_454/merge_stmt_1735_PhiAck/$entry
      -- CP-element group 269: 	 branch_block_stmt_454/merge_stmt_1735_PhiAck/$exit
      -- CP-element group 269: 	 branch_block_stmt_454/merge_stmt_1735_PhiReqMerge
      -- CP-element group 269: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/$exit
      -- CP-element group 269: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_454/call_stmt_1719_to_assign_stmt_1732/WPIPE_elapsed_time_pipe_1730_Update/ack
      -- CP-element group 269: 	 branch_block_stmt_454/return___PhiReq/$entry
      -- CP-element group 269: 	 branch_block_stmt_454/return___PhiReq/$exit
      -- CP-element group 269: 	 branch_block_stmt_454/merge_stmt_1735_PhiAck/dummy
      -- 
    ack_3308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1730_inst_ack_1, ack => convolution3D_CP_1129_elements(269)); -- 
    -- CP-element group 270:  transition  output  delay-element  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	86 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	274 
    -- CP-element group 270:  members (5) 
      -- CP-element group 270: 	 branch_block_stmt_454/bbx_xnph327_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_req
      -- CP-element group 270: 	 branch_block_stmt_454/bbx_xnph327_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770_konst_delay_trans
      -- CP-element group 270: 	 branch_block_stmt_454/bbx_xnph327_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/$exit
      -- CP-element group 270: 	 branch_block_stmt_454/bbx_xnph327_forx_xbody_PhiReq/phi_stmt_764/$exit
      -- CP-element group 270: 	 branch_block_stmt_454/bbx_xnph327_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_764_req_3331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_764_req_3331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(270), ack => phi_stmt_764_req_1); -- 
    -- Element group convolution3D_CP_1129_elements(270) is a control-delay.
    cp_element_270_delay: control_delay_element  generic map(name => " 270_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(86), ack => convolution3D_CP_1129_elements(270), clk => clk, reset =>reset);
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	128 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	273 
    -- CP-element group 271:  members (2) 
      -- CP-element group 271: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/SplitProtocol/Sample/ra
      -- CP-element group 271: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/SplitProtocol/Sample/$exit
      -- 
    ra_3351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_767_inst_ack_0, ack => convolution3D_CP_1129_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	128 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (2) 
      -- CP-element group 272: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/SplitProtocol/Update/ca
      -- CP-element group 272: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/SplitProtocol/Update/$exit
      -- 
    ca_3356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_767_inst_ack_1, ack => convolution3D_CP_1129_elements(272)); -- 
    -- CP-element group 273:  join  transition  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/$exit
      -- CP-element group 273: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_req
      -- CP-element group 273: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/SplitProtocol/$exit
      -- CP-element group 273: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_767/$exit
      -- CP-element group 273: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 273: 	 branch_block_stmt_454/forx_xbody_forx_xbody_PhiReq/phi_stmt_764/phi_stmt_764_sources/$exit
      -- 
    phi_stmt_764_req_3357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_764_req_3357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(273), ack => phi_stmt_764_req_0); -- 
    convolution3D_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(271) & convolution3D_CP_1129_elements(272);
      gj_convolution3D_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  merge  transition  place  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	270 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_454/merge_stmt_763_PhiAck/$entry
      -- CP-element group 274: 	 branch_block_stmt_454/merge_stmt_763_PhiReqMerge
      -- 
    convolution3D_CP_1129_elements(274) <= OrReduce(convolution3D_CP_1129_elements(270) & convolution3D_CP_1129_elements(273));
    -- CP-element group 275:  fork  transition  place  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	87 
    -- CP-element group 275: 	88 
    -- CP-element group 275: 	90 
    -- CP-element group 275: 	91 
    -- CP-element group 275: 	94 
    -- CP-element group 275: 	98 
    -- CP-element group 275: 	102 
    -- CP-element group 275: 	106 
    -- CP-element group 275: 	110 
    -- CP-element group 275: 	114 
    -- CP-element group 275: 	118 
    -- CP-element group 275: 	122 
    -- CP-element group 275: 	125 
    -- CP-element group 275:  members (56) 
      -- CP-element group 275: 	 branch_block_stmt_454/merge_stmt_763__exit__
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926__entry__
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_update_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_resized_1
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_scaled_1
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_computed_1
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_resize_1/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_resize_1/$exit
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_resize_1/index_resize_req
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_resize_1/index_resize_ack
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_scale_1/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_scale_1/$exit
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_scale_1/scale_rename_req
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_scale_1/scale_rename_ack
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_update_start
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Sample/req
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Update/req
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_complete/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/addr_of_777_complete/req
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/RPIPE_maxpool_input_pipe_780_Sample/rr
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_update_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_784_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_update_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_797_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_update_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_815_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_update_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_833_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_update_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_851_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_update_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_869_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_update_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_887_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_update_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/type_cast_905_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_update_start_
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/word_0/$entry
      -- CP-element group 275: 	 branch_block_stmt_454/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/word_0/cr
      -- CP-element group 275: 	 branch_block_stmt_454/merge_stmt_763_PhiAck/phi_stmt_764_ack
      -- CP-element group 275: 	 branch_block_stmt_454/merge_stmt_763_PhiAck/$exit
      -- 
    phi_stmt_764_ack_3362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_764_ack_0, ack => convolution3D_CP_1129_elements(275)); -- 
    req_1833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => array_obj_ref_776_index_offset_req_0); -- 
    req_1838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => array_obj_ref_776_index_offset_req_1); -- 
    req_1853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => addr_of_777_final_reg_req_1); -- 
    rr_1862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => RPIPE_maxpool_input_pipe_780_inst_req_0); -- 
    cr_1881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => type_cast_784_inst_req_1); -- 
    cr_1909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => type_cast_797_inst_req_1); -- 
    cr_1937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => type_cast_815_inst_req_1); -- 
    cr_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => type_cast_833_inst_req_1); -- 
    cr_1993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => type_cast_851_inst_req_1); -- 
    cr_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => type_cast_869_inst_req_1); -- 
    cr_2049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => type_cast_887_inst_req_1); -- 
    cr_2077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => type_cast_905_inst_req_1); -- 
    cr_2127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(275), ack => ptr_deref_913_store_0_req_1); -- 
    -- CP-element group 276:  transition  output  delay-element  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	76 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	280 
    -- CP-element group 276:  members (5) 
      -- CP-element group 276: 	 branch_block_stmt_454/entry_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/$exit
      -- CP-element group 276: 	 branch_block_stmt_454/entry_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_964_konst_delay_trans
      -- CP-element group 276: 	 branch_block_stmt_454/entry_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_req
      -- CP-element group 276: 	 branch_block_stmt_454/entry_forx_xend_PhiReq/phi_stmt_958/$exit
      -- CP-element group 276: 	 branch_block_stmt_454/entry_forx_xend_PhiReq/$exit
      -- 
    phi_stmt_958_req_3385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_958_req_3385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(276), ack => phi_stmt_958_req_1); -- 
    -- Element group convolution3D_CP_1129_elements(276) is a control-delay.
    cp_element_276_delay: control_delay_element  generic map(name => " 276_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(76), ack => convolution3D_CP_1129_elements(276), clk => clk, reset =>reset);
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	127 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (2) 
      -- CP-element group 277: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/SplitProtocol/Sample/ra
      -- CP-element group 277: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/SplitProtocol/Sample/$exit
      -- 
    ra_3405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_961_inst_ack_0, ack => convolution3D_CP_1129_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	127 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (2) 
      -- CP-element group 278: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/SplitProtocol/Update/ca
      -- CP-element group 278: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/SplitProtocol/Update/$exit
      -- 
    ca_3410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_961_inst_ack_1, ack => convolution3D_CP_1129_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/$exit
      -- CP-element group 279: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/$exit
      -- CP-element group 279: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_req
      -- CP-element group 279: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 279: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/SplitProtocol/$exit
      -- CP-element group 279: 	 branch_block_stmt_454/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_958/phi_stmt_958_sources/type_cast_961/$exit
      -- 
    phi_stmt_958_req_3411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_958_req_3411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(279), ack => phi_stmt_958_req_0); -- 
    convolution3D_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(277) & convolution3D_CP_1129_elements(278);
      gj_convolution3D_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  merge  transition  place  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	276 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (2) 
      -- CP-element group 280: 	 branch_block_stmt_454/merge_stmt_957_PhiReqMerge
      -- CP-element group 280: 	 branch_block_stmt_454/merge_stmt_957_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(280) <= OrReduce(convolution3D_CP_1129_elements(276) & convolution3D_CP_1129_elements(279));
    -- CP-element group 281:  branch  transition  place  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	129 
    -- CP-element group 281: 	130 
    -- CP-element group 281:  members (15) 
      -- CP-element group 281: 	 branch_block_stmt_454/merge_stmt_957__exit__
      -- CP-element group 281: 	 branch_block_stmt_454/assign_stmt_971_to_assign_stmt_977__entry__
      -- CP-element group 281: 	 branch_block_stmt_454/assign_stmt_971_to_assign_stmt_977__exit__
      -- CP-element group 281: 	 branch_block_stmt_454/if_stmt_978__entry__
      -- CP-element group 281: 	 branch_block_stmt_454/assign_stmt_971_to_assign_stmt_977/$entry
      -- CP-element group 281: 	 branch_block_stmt_454/assign_stmt_971_to_assign_stmt_977/$exit
      -- CP-element group 281: 	 branch_block_stmt_454/if_stmt_978_dead_link/$entry
      -- CP-element group 281: 	 branch_block_stmt_454/if_stmt_978_eval_test/$entry
      -- CP-element group 281: 	 branch_block_stmt_454/if_stmt_978_eval_test/$exit
      -- CP-element group 281: 	 branch_block_stmt_454/if_stmt_978_eval_test/branch_req
      -- CP-element group 281: 	 branch_block_stmt_454/R_tobool_979_place
      -- CP-element group 281: 	 branch_block_stmt_454/if_stmt_978_if_link/$entry
      -- CP-element group 281: 	 branch_block_stmt_454/if_stmt_978_else_link/$entry
      -- CP-element group 281: 	 branch_block_stmt_454/merge_stmt_957_PhiAck/phi_stmt_958_ack
      -- CP-element group 281: 	 branch_block_stmt_454/merge_stmt_957_PhiAck/$exit
      -- 
    phi_stmt_958_ack_3416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_958_ack_0, ack => convolution3D_CP_1129_elements(281)); -- 
    branch_req_2161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(281), ack => if_stmt_978_branch_req_0); -- 
    -- CP-element group 282:  transition  output  delay-element  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	130 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (4) 
      -- CP-element group 282: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_req
      -- CP-element group 282: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1003_konst_delay_trans
      -- CP-element group 282: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/$exit
      -- CP-element group 282: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/$exit
      -- 
    phi_stmt_999_req_3439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_999_req_3439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(282), ack => phi_stmt_999_req_0); -- 
    -- Element group convolution3D_CP_1129_elements(282) is a control-delay.
    cp_element_282_delay: control_delay_element  generic map(name => " 282_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(130), ack => convolution3D_CP_1129_elements(282), clk => clk, reset =>reset);
    -- CP-element group 283:  transition  output  delay-element  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	130 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (4) 
      -- CP-element group 283: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_req
      -- CP-element group 283: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1010_konst_delay_trans
      -- CP-element group 283: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/$exit
      -- CP-element group 283: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/$exit
      -- 
    phi_stmt_1006_req_3447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1006_req_3447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(283), ack => phi_stmt_1006_req_0); -- 
    -- Element group convolution3D_CP_1129_elements(283) is a control-delay.
    cp_element_283_delay: control_delay_element  generic map(name => " 283_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(130), ack => convolution3D_CP_1129_elements(283), clk => clk, reset =>reset);
    -- CP-element group 284:  join  transition  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	292 
    -- CP-element group 284:  members (1) 
      -- CP-element group 284: 	 branch_block_stmt_454/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(282) & convolution3D_CP_1129_elements(283);
      gj_convolution3D_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	138 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (2) 
      -- CP-element group 285: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Sample/ra
      -- CP-element group 285: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Sample/$exit
      -- 
    ra_3467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_0, ack => convolution3D_CP_1129_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	138 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Update/ca
      -- 
    ca_3472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_1, ack => convolution3D_CP_1129_elements(286)); -- 
    -- CP-element group 287:  join  transition  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	291 
    -- CP-element group 287:  members (5) 
      -- CP-element group 287: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_req
      -- CP-element group 287: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/$exit
      -- CP-element group 287: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/$exit
      -- CP-element group 287: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/phi_stmt_999_sources/$exit
      -- CP-element group 287: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_999/$exit
      -- 
    phi_stmt_999_req_3473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_999_req_3473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(287), ack => phi_stmt_999_req_1); -- 
    convolution3D_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(285) & convolution3D_CP_1129_elements(286);
      gj_convolution3D_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  transition  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	138 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (2) 
      -- CP-element group 288: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/SplitProtocol/Sample/ra
      -- CP-element group 288: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/SplitProtocol/Sample/$exit
      -- 
    ra_3490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1012_inst_ack_0, ack => convolution3D_CP_1129_elements(288)); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	138 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (2) 
      -- CP-element group 289: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/SplitProtocol/Update/ca
      -- CP-element group 289: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/SplitProtocol/Update/$exit
      -- 
    ca_3495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1012_inst_ack_1, ack => convolution3D_CP_1129_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (5) 
      -- CP-element group 290: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_req
      -- CP-element group 290: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/SplitProtocol/$exit
      -- CP-element group 290: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/type_cast_1012/$exit
      -- CP-element group 290: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/phi_stmt_1006_sources/$exit
      -- CP-element group 290: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1006/$exit
      -- 
    phi_stmt_1006_req_3496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1006_req_3496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(290), ack => phi_stmt_1006_req_1); -- 
    convolution3D_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(288) & convolution3D_CP_1129_elements(289);
      gj_convolution3D_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  join  transition  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	287 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (1) 
      -- CP-element group 291: 	 branch_block_stmt_454/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(287) & convolution3D_CP_1129_elements(290);
      gj_convolution3D_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  merge  fork  transition  place  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	284 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292: 	294 
    -- CP-element group 292:  members (2) 
      -- CP-element group 292: 	 branch_block_stmt_454/merge_stmt_998_PhiReqMerge
      -- CP-element group 292: 	 branch_block_stmt_454/merge_stmt_998_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(292) <= OrReduce(convolution3D_CP_1129_elements(284) & convolution3D_CP_1129_elements(291));
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (1) 
      -- CP-element group 293: 	 branch_block_stmt_454/merge_stmt_998_PhiAck/phi_stmt_999_ack
      -- 
    phi_stmt_999_ack_3501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_999_ack_0, ack => convolution3D_CP_1129_elements(293)); -- 
    -- CP-element group 294:  transition  input  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	292 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (1) 
      -- CP-element group 294: 	 branch_block_stmt_454/merge_stmt_998_PhiAck/phi_stmt_1006_ack
      -- 
    phi_stmt_1006_ack_3502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1006_ack_0, ack => convolution3D_CP_1129_elements(294)); -- 
    -- CP-element group 295:  join  fork  transition  place  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	131 
    -- CP-element group 295: 	134 
    -- CP-element group 295: 	135 
    -- CP-element group 295: 	136 
    -- CP-element group 295:  members (16) 
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_update_start_
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_Sample/rr
      -- CP-element group 295: 	 branch_block_stmt_454/merge_stmt_998__exit__
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052__entry__
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_sample_start_
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1046_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/$entry
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_sample_start_
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/RPIPE_maxpool_input_pipe_1027_Sample/rr
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_update_start_
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_454/assign_stmt_1019_to_assign_stmt_1052/type_cast_1031_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_454/merge_stmt_998_PhiAck/$exit
      -- 
    rr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(295), ack => type_cast_1046_inst_req_0); -- 
    cr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(295), ack => type_cast_1046_inst_req_1); -- 
    rr_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(295), ack => RPIPE_maxpool_input_pipe_1027_inst_req_0); -- 
    cr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(295), ack => type_cast_1031_inst_req_1); -- 
    convolution3D_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(293) & convolution3D_CP_1129_elements(294);
      gj_convolution3D_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	139 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	298 
    -- CP-element group 296:  members (2) 
      -- CP-element group 296: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/SplitProtocol/Sample/ra
      -- CP-element group 296: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/SplitProtocol/Sample/$exit
      -- 
    ra_3526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1063_inst_ack_0, ack => convolution3D_CP_1129_elements(296)); -- 
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	139 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (2) 
      -- CP-element group 297: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/SplitProtocol/Update/ca
      -- CP-element group 297: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/SplitProtocol/Update/$exit
      -- 
    ca_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1063_inst_ack_1, ack => convolution3D_CP_1129_elements(297)); -- 
    -- CP-element group 298:  join  transition  place  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	296 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (8) 
      -- CP-element group 298: 	 branch_block_stmt_454/merge_stmt_1059_PhiReqMerge
      -- CP-element group 298: 	 branch_block_stmt_454/merge_stmt_1059_PhiAck/$entry
      -- CP-element group 298: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_req
      -- CP-element group 298: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/SplitProtocol/$exit
      -- CP-element group 298: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/type_cast_1063/$exit
      -- CP-element group 298: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/phi_stmt_1060_sources/$exit
      -- CP-element group 298: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1060/$exit
      -- CP-element group 298: 	 branch_block_stmt_454/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- 
    phi_stmt_1060_req_3532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1060_req_3532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(298), ack => phi_stmt_1060_req_0); -- 
    convolution3D_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(296) & convolution3D_CP_1129_elements(297);
      gj_convolution3D_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	140 
    -- CP-element group 299: 	141 
    -- CP-element group 299: 	143 
    -- CP-element group 299: 	145 
    -- CP-element group 299:  members (29) 
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_scale_1/scale_rename_ack
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_final_index_sum_regn_update_start
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_final_index_sum_regn_Sample/$entry
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Update/word_access_complete/$entry
      -- CP-element group 299: 	 branch_block_stmt_454/merge_stmt_1059__exit__
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098__entry__
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/$entry
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_update_start_
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_scale_1/scale_rename_req
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_scale_1/$exit
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_scale_1/$entry
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_resize_1/index_resize_ack
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_resize_1/index_resize_req
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_resize_1/$exit
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_resize_1/$entry
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_computed_1
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_scaled_1
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_index_resized_1
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_update_start_
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_final_index_sum_regn_Update/req
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_final_index_sum_regn_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_complete/req
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Update/word_access_complete/word_0/cr
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/addr_of_1093_complete/$entry
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/ptr_deref_1096_Update/word_access_complete/word_0/$entry
      -- CP-element group 299: 	 branch_block_stmt_454/assign_stmt_1070_to_assign_stmt_1098/array_obj_ref_1092_final_index_sum_regn_Sample/req
      -- CP-element group 299: 	 branch_block_stmt_454/merge_stmt_1059_PhiAck/phi_stmt_1060_ack
      -- CP-element group 299: 	 branch_block_stmt_454/merge_stmt_1059_PhiAck/$exit
      -- 
    phi_stmt_1060_ack_3537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1060_ack_0, ack => convolution3D_CP_1129_elements(299)); -- 
    req_2272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(299), ack => array_obj_ref_1092_index_offset_req_1); -- 
    req_2287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(299), ack => addr_of_1093_final_reg_req_1); -- 
    cr_2337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(299), ack => ptr_deref_1096_store_0_req_1); -- 
    req_2267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(299), ack => array_obj_ref_1092_index_offset_req_0); -- 
    -- CP-element group 300:  merge  fork  transition  place  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	129 
    -- CP-element group 300: 	146 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	147 
    -- CP-element group 300: 	148 
    -- CP-element group 300: 	149 
    -- CP-element group 300: 	150 
    -- CP-element group 300: 	151 
    -- CP-element group 300: 	152 
    -- CP-element group 300: 	153 
    -- CP-element group 300: 	154 
    -- CP-element group 300:  members (31) 
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_Sample/rr
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_Update/cr
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_454/merge_stmt_1100__exit__
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152__entry__
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_update_start_
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_Update/cr
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_Sample/rr
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_update_start_
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1115_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_Update/cr
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_454/merge_stmt_1100_PhiReqMerge
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_Sample/rr
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_update_start_
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1111_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_Update/cr
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_Sample/rr
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1103_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/$entry
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_454/assign_stmt_1104_to_assign_stmt_1152/type_cast_1107_update_start_
      -- CP-element group 300: 	 branch_block_stmt_454/merge_stmt_1100_PhiAck/dummy
      -- CP-element group 300: 	 branch_block_stmt_454/merge_stmt_1100_PhiAck/$exit
      -- CP-element group 300: 	 branch_block_stmt_454/merge_stmt_1100_PhiAck/$entry
      -- 
    rr_2349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(300), ack => type_cast_1103_inst_req_0); -- 
    cr_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(300), ack => type_cast_1103_inst_req_1); -- 
    cr_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(300), ack => type_cast_1115_inst_req_1); -- 
    rr_2391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(300), ack => type_cast_1115_inst_req_0); -- 
    cr_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(300), ack => type_cast_1111_inst_req_1); -- 
    rr_2377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(300), ack => type_cast_1111_inst_req_0); -- 
    cr_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(300), ack => type_cast_1107_inst_req_1); -- 
    rr_2363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(300), ack => type_cast_1107_inst_req_0); -- 
    convolution3D_CP_1129_elements(300) <= OrReduce(convolution3D_CP_1129_elements(129) & convolution3D_CP_1129_elements(146));
    -- CP-element group 301:  transition  output  delay-element  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	170 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	305 
    -- CP-element group 301:  members (5) 
      -- CP-element group 301: 	 branch_block_stmt_454/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_req
      -- CP-element group 301: 	 branch_block_stmt_454/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1237_konst_delay_trans
      -- CP-element group 301: 	 branch_block_stmt_454/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/$exit
      -- CP-element group 301: 	 branch_block_stmt_454/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1233/$exit
      -- CP-element group 301: 	 branch_block_stmt_454/bbx_xnph_forx_xbody163_PhiReq/$exit
      -- 
    phi_stmt_1233_req_3571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1233_req_3571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(301), ack => phi_stmt_1233_req_0); -- 
    -- Element group convolution3D_CP_1129_elements(301) is a control-delay.
    cp_element_301_delay: control_delay_element  generic map(name => " 301_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(170), ack => convolution3D_CP_1129_elements(301), clk => clk, reset =>reset);
    -- CP-element group 302:  transition  input  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	212 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (2) 
      -- CP-element group 302: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/SplitProtocol/Sample/ra
      -- CP-element group 302: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/SplitProtocol/Sample/$exit
      -- 
    ra_3591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1239_inst_ack_0, ack => convolution3D_CP_1129_elements(302)); -- 
    -- CP-element group 303:  transition  input  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	212 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (2) 
      -- CP-element group 303: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/SplitProtocol/Update/$exit
      -- CP-element group 303: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/SplitProtocol/Update/ca
      -- 
    ca_3596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1239_inst_ack_1, ack => convolution3D_CP_1129_elements(303)); -- 
    -- CP-element group 304:  join  transition  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/SplitProtocol/$exit
      -- CP-element group 304: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/type_cast_1239/$exit
      -- CP-element group 304: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_sources/$exit
      -- CP-element group 304: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/$exit
      -- CP-element group 304: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/$exit
      -- CP-element group 304: 	 branch_block_stmt_454/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1233/phi_stmt_1233_req
      -- 
    phi_stmt_1233_req_3597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1233_req_3597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(304), ack => phi_stmt_1233_req_1); -- 
    convolution3D_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(302) & convolution3D_CP_1129_elements(303);
      gj_convolution3D_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  merge  transition  place  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	301 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (2) 
      -- CP-element group 305: 	 branch_block_stmt_454/merge_stmt_1232_PhiReqMerge
      -- CP-element group 305: 	 branch_block_stmt_454/merge_stmt_1232_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(305) <= OrReduce(convolution3D_CP_1129_elements(301) & convolution3D_CP_1129_elements(304));
    -- CP-element group 306:  fork  transition  place  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	171 
    -- CP-element group 306: 	172 
    -- CP-element group 306: 	174 
    -- CP-element group 306: 	175 
    -- CP-element group 306: 	178 
    -- CP-element group 306: 	182 
    -- CP-element group 306: 	186 
    -- CP-element group 306: 	190 
    -- CP-element group 306: 	194 
    -- CP-element group 306: 	198 
    -- CP-element group 306: 	202 
    -- CP-element group 306: 	206 
    -- CP-element group 306: 	209 
    -- CP-element group 306:  members (56) 
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_Update/cr
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_final_index_sum_regn_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_final_index_sum_regn_update_start
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_final_index_sum_regn_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_final_index_sum_regn_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_update_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_final_index_sum_regn_Update/req
      -- CP-element group 306: 	 branch_block_stmt_454/merge_stmt_1232__exit__
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395__entry__
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_Update/cr
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_scale_1/scale_rename_ack
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_scale_1/scale_rename_req
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_scale_1/$exit
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_scale_1/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_resize_1/index_resize_ack
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_resize_1/index_resize_req
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_update_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_resize_1/$exit
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_resize_1/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_update_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_computed_1
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_scaled_1
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/array_obj_ref_1245_index_resized_1
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1253_update_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_Update/cr
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_update_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1266_update_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_Sample/rr
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_Update/cr
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1320_Update/cr
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_complete/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1284_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1302_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/RPIPE_maxpool_input_pipe_1249_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/addr_of_1246_complete/req
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_update_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1338_Update/cr
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_update_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1356_Update/cr
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_update_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/type_cast_1374_Update/cr
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_update_start_
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Update/word_access_complete/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Update/word_access_complete/word_0/$entry
      -- CP-element group 306: 	 branch_block_stmt_454/assign_stmt_1247_to_assign_stmt_1395/ptr_deref_1382_Update/word_access_complete/word_0/cr
      -- CP-element group 306: 	 branch_block_stmt_454/merge_stmt_1232_PhiAck/phi_stmt_1233_ack
      -- CP-element group 306: 	 branch_block_stmt_454/merge_stmt_1232_PhiAck/$exit
      -- 
    phi_stmt_1233_ack_3602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1233_ack_0, ack => convolution3D_CP_1129_elements(306)); -- 
    cr_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => type_cast_1302_inst_req_1); -- 
    req_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => array_obj_ref_1245_index_offset_req_0); -- 
    req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => array_obj_ref_1245_index_offset_req_1); -- 
    cr_2579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => type_cast_1253_inst_req_1); -- 
    cr_2607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => type_cast_1266_inst_req_1); -- 
    rr_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => RPIPE_maxpool_input_pipe_1249_inst_req_0); -- 
    cr_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => type_cast_1284_inst_req_1); -- 
    cr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => type_cast_1320_inst_req_1); -- 
    req_2551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => addr_of_1246_final_reg_req_1); -- 
    cr_2719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => type_cast_1338_inst_req_1); -- 
    cr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => type_cast_1356_inst_req_1); -- 
    cr_2775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => type_cast_1374_inst_req_1); -- 
    cr_2825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(306), ack => ptr_deref_1382_store_0_req_1); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	211 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	309 
    -- CP-element group 307:  members (2) 
      -- CP-element group 307: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Sample/ra
      -- CP-element group 307: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Sample/$exit
      -- 
    ra_3634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1430_inst_ack_0, ack => convolution3D_CP_1129_elements(307)); -- 
    -- CP-element group 308:  transition  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	211 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (2) 
      -- CP-element group 308: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Update/ca
      -- CP-element group 308: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/Update/$exit
      -- 
    ca_3639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1430_inst_ack_1, ack => convolution3D_CP_1129_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	307 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$exit
      -- CP-element group 309: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_req
      -- CP-element group 309: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/$exit
      -- CP-element group 309: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$exit
      -- CP-element group 309: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/SplitProtocol/$exit
      -- CP-element group 309: 	 branch_block_stmt_454/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1430/$exit
      -- 
    phi_stmt_1427_req_3640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1427_req_3640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(309), ack => phi_stmt_1427_req_0); -- 
    convolution3D_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(307) & convolution3D_CP_1129_elements(308);
      gj_convolution3D_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  transition  output  delay-element  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	157 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (5) 
      -- CP-element group 310: 	 branch_block_stmt_454/ifx_xend_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_req
      -- CP-element group 310: 	 branch_block_stmt_454/ifx_xend_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/type_cast_1433_konst_delay_trans
      -- CP-element group 310: 	 branch_block_stmt_454/ifx_xend_forx_xend215_PhiReq/phi_stmt_1427/phi_stmt_1427_sources/$exit
      -- CP-element group 310: 	 branch_block_stmt_454/ifx_xend_forx_xend215_PhiReq/phi_stmt_1427/$exit
      -- CP-element group 310: 	 branch_block_stmt_454/ifx_xend_forx_xend215_PhiReq/$exit
      -- 
    phi_stmt_1427_req_3651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1427_req_3651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(310), ack => phi_stmt_1427_req_1); -- 
    -- Element group convolution3D_CP_1129_elements(310) is a control-delay.
    cp_element_310_delay: control_delay_element  generic map(name => " 310_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(157), ack => convolution3D_CP_1129_elements(310), clk => clk, reset =>reset);
    -- CP-element group 311:  merge  transition  place  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (2) 
      -- CP-element group 311: 	 branch_block_stmt_454/merge_stmt_1426_PhiReqMerge
      -- CP-element group 311: 	 branch_block_stmt_454/merge_stmt_1426_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(311) <= OrReduce(convolution3D_CP_1129_elements(309) & convolution3D_CP_1129_elements(310));
    -- CP-element group 312:  branch  transition  place  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	213 
    -- CP-element group 312: 	214 
    -- CP-element group 312:  members (15) 
      -- CP-element group 312: 	 branch_block_stmt_454/merge_stmt_1426_PhiAck/phi_stmt_1427_ack
      -- CP-element group 312: 	 branch_block_stmt_454/merge_stmt_1426__exit__
      -- CP-element group 312: 	 branch_block_stmt_454/assign_stmt_1440_to_assign_stmt_1446__entry__
      -- CP-element group 312: 	 branch_block_stmt_454/assign_stmt_1440_to_assign_stmt_1446__exit__
      -- CP-element group 312: 	 branch_block_stmt_454/if_stmt_1447__entry__
      -- CP-element group 312: 	 branch_block_stmt_454/merge_stmt_1426_PhiAck/$exit
      -- CP-element group 312: 	 branch_block_stmt_454/assign_stmt_1440_to_assign_stmt_1446/$entry
      -- CP-element group 312: 	 branch_block_stmt_454/assign_stmt_1440_to_assign_stmt_1446/$exit
      -- CP-element group 312: 	 branch_block_stmt_454/if_stmt_1447_dead_link/$entry
      -- CP-element group 312: 	 branch_block_stmt_454/if_stmt_1447_eval_test/$entry
      -- CP-element group 312: 	 branch_block_stmt_454/if_stmt_1447_eval_test/$exit
      -- CP-element group 312: 	 branch_block_stmt_454/if_stmt_1447_eval_test/branch_req
      -- CP-element group 312: 	 branch_block_stmt_454/R_tobool218_1448_place
      -- CP-element group 312: 	 branch_block_stmt_454/if_stmt_1447_if_link/$entry
      -- CP-element group 312: 	 branch_block_stmt_454/if_stmt_1447_else_link/$entry
      -- 
    phi_stmt_1427_ack_3656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1427_ack_0, ack => convolution3D_CP_1129_elements(312)); -- 
    branch_req_2859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => if_stmt_1447_branch_req_0); -- 
    -- CP-element group 313:  transition  output  delay-element  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	216 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	315 
    -- CP-element group 313:  members (4) 
      -- CP-element group 313: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_req
      -- CP-element group 313: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1476_konst_delay_trans
      -- CP-element group 313: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/$exit
      -- CP-element group 313: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/$exit
      -- 
    phi_stmt_1472_req_3679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1472_req_3679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(313), ack => phi_stmt_1472_req_0); -- 
    -- Element group convolution3D_CP_1129_elements(313) is a control-delay.
    cp_element_313_delay: control_delay_element  generic map(name => " 313_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(216), ack => convolution3D_CP_1129_elements(313), clk => clk, reset =>reset);
    -- CP-element group 314:  transition  output  delay-element  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	216 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (4) 
      -- CP-element group 314: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_req
      -- CP-element group 314: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1483_konst_delay_trans
      -- CP-element group 314: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/$exit
      -- CP-element group 314: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/$exit
      -- 
    phi_stmt_1479_req_3687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1479_req_3687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(314), ack => phi_stmt_1479_req_0); -- 
    -- Element group convolution3D_CP_1129_elements(314) is a control-delay.
    cp_element_314_delay: control_delay_element  generic map(name => " 314_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(216), ack => convolution3D_CP_1129_elements(314), clk => clk, reset =>reset);
    -- CP-element group 315:  join  transition  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	313 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	323 
    -- CP-element group 315:  members (1) 
      -- CP-element group 315: 	 branch_block_stmt_454/bbx_xnphx_xi298_forx_xbodyx_xi307_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(313) & convolution3D_CP_1129_elements(314);
      gj_convolution3D_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	224 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	318 
    -- CP-element group 316:  members (2) 
      -- CP-element group 316: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/SplitProtocol/Sample/ra
      -- CP-element group 316: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/SplitProtocol/Sample/$exit
      -- 
    ra_3707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1478_inst_ack_0, ack => convolution3D_CP_1129_elements(316)); -- 
    -- CP-element group 317:  transition  input  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	224 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (2) 
      -- CP-element group 317: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/SplitProtocol/Update/ca
      -- CP-element group 317: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/SplitProtocol/Update/$exit
      -- 
    ca_3712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1478_inst_ack_1, ack => convolution3D_CP_1129_elements(317)); -- 
    -- CP-element group 318:  join  transition  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	316 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	322 
    -- CP-element group 318:  members (5) 
      -- CP-element group 318: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/SplitProtocol/$exit
      -- CP-element group 318: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/type_cast_1478/$exit
      -- CP-element group 318: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_sources/$exit
      -- CP-element group 318: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/$exit
      -- CP-element group 318: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1472/phi_stmt_1472_req
      -- 
    phi_stmt_1472_req_3713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1472_req_3713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(318), ack => phi_stmt_1472_req_1); -- 
    convolution3D_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(316) & convolution3D_CP_1129_elements(317);
      gj_convolution3D_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	224 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (2) 
      -- CP-element group 319: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/SplitProtocol/Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/SplitProtocol/Sample/ra
      -- 
    ra_3730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1485_inst_ack_0, ack => convolution3D_CP_1129_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	224 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (2) 
      -- CP-element group 320: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/SplitProtocol/Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/SplitProtocol/Update/ca
      -- 
    ca_3735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1485_inst_ack_1, ack => convolution3D_CP_1129_elements(320)); -- 
    -- CP-element group 321:  join  transition  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (5) 
      -- CP-element group 321: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/$exit
      -- CP-element group 321: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/type_cast_1485/SplitProtocol/$exit
      -- CP-element group 321: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_sources/$exit
      -- CP-element group 321: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/$exit
      -- CP-element group 321: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/phi_stmt_1479/phi_stmt_1479_req
      -- 
    phi_stmt_1479_req_3736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1479_req_3736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(321), ack => phi_stmt_1479_req_1); -- 
    convolution3D_cp_element_group_321: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_321"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(319) & convolution3D_CP_1129_elements(320);
      gj_convolution3D_cp_element_group_321 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(321), clk => clk, reset => reset); --
    end block;
    -- CP-element group 322:  join  transition  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	318 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (1) 
      -- CP-element group 322: 	 branch_block_stmt_454/forx_xbodyx_xi307_forx_xbodyx_xi307_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(318) & convolution3D_CP_1129_elements(321);
      gj_convolution3D_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  merge  fork  transition  place  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	315 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (2) 
      -- CP-element group 323: 	 branch_block_stmt_454/merge_stmt_1471_PhiReqMerge
      -- CP-element group 323: 	 branch_block_stmt_454/merge_stmt_1471_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(323) <= OrReduce(convolution3D_CP_1129_elements(315) & convolution3D_CP_1129_elements(322));
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (1) 
      -- CP-element group 324: 	 branch_block_stmt_454/merge_stmt_1471_PhiAck/phi_stmt_1472_ack
      -- 
    phi_stmt_1472_ack_3741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1472_ack_0, ack => convolution3D_CP_1129_elements(324)); -- 
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (1) 
      -- CP-element group 325: 	 branch_block_stmt_454/merge_stmt_1471_PhiAck/phi_stmt_1479_ack
      -- 
    phi_stmt_1479_ack_3742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1479_ack_0, ack => convolution3D_CP_1129_elements(325)); -- 
    -- CP-element group 326:  join  fork  transition  place  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	217 
    -- CP-element group 326: 	220 
    -- CP-element group 326: 	221 
    -- CP-element group 326: 	222 
    -- CP-element group 326:  members (16) 
      -- CP-element group 326: 	 branch_block_stmt_454/merge_stmt_1471__exit__
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525__entry__
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/$entry
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/RPIPE_maxpool_input_pipe_1500_Sample/rr
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_update_start_
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1504_Update/cr
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_update_start_
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_Sample/rr
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_454/assign_stmt_1492_to_assign_stmt_1525/type_cast_1519_Update/cr
      -- CP-element group 326: 	 branch_block_stmt_454/merge_stmt_1471_PhiAck/$exit
      -- 
    rr_2898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(326), ack => RPIPE_maxpool_input_pipe_1500_inst_req_0); -- 
    cr_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(326), ack => type_cast_1504_inst_req_1); -- 
    rr_2926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(326), ack => type_cast_1519_inst_req_0); -- 
    cr_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(326), ack => type_cast_1519_inst_req_1); -- 
    convolution3D_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(324) & convolution3D_CP_1129_elements(325);
      gj_convolution3D_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	225 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	329 
    -- CP-element group 327:  members (2) 
      -- CP-element group 327: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/SplitProtocol/Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/SplitProtocol/Sample/ra
      -- 
    ra_3766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1536_inst_ack_0, ack => convolution3D_CP_1129_elements(327)); -- 
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	225 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (2) 
      -- CP-element group 328: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/SplitProtocol/Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/SplitProtocol/Update/ca
      -- 
    ca_3771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1536_inst_ack_1, ack => convolution3D_CP_1129_elements(328)); -- 
    -- CP-element group 329:  join  transition  place  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	327 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (8) 
      -- CP-element group 329: 	 branch_block_stmt_454/merge_stmt_1532_PhiReqMerge
      -- CP-element group 329: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/$exit
      -- CP-element group 329: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/$exit
      -- CP-element group 329: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/$exit
      -- CP-element group 329: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/$exit
      -- CP-element group 329: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_sources/type_cast_1536/SplitProtocol/$exit
      -- CP-element group 329: 	 branch_block_stmt_454/forx_xbodyx_xi307_getRemainingElementsx_xexit315_PhiReq/phi_stmt_1533/phi_stmt_1533_req
      -- CP-element group 329: 	 branch_block_stmt_454/merge_stmt_1532_PhiAck/$entry
      -- 
    phi_stmt_1533_req_3772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1533_req_3772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(329), ack => phi_stmt_1533_req_0); -- 
    convolution3D_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(327) & convolution3D_CP_1129_elements(328);
      gj_convolution3D_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	226 
    -- CP-element group 330: 	227 
    -- CP-element group 330: 	229 
    -- CP-element group 330: 	231 
    -- CP-element group 330:  members (29) 
      -- CP-element group 330: 	 branch_block_stmt_454/merge_stmt_1532__exit__
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571__entry__
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/$entry
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_update_start_
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_resized_1
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_scaled_1
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_computed_1
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_resize_1/$entry
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_resize_1/$exit
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_resize_1/index_resize_req
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_resize_1/index_resize_ack
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_scale_1/$entry
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_scale_1/$exit
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_scale_1/scale_rename_req
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_index_scale_1/scale_rename_ack
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_final_index_sum_regn_update_start
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_final_index_sum_regn_Sample/$entry
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_final_index_sum_regn_Sample/req
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_final_index_sum_regn_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/array_obj_ref_1565_final_index_sum_regn_Update/req
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_complete/$entry
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/addr_of_1566_complete/req
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_update_start_
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Update/word_access_complete/$entry
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Update/word_access_complete/word_0/$entry
      -- CP-element group 330: 	 branch_block_stmt_454/assign_stmt_1543_to_assign_stmt_1571/ptr_deref_1569_Update/word_access_complete/word_0/cr
      -- CP-element group 330: 	 branch_block_stmt_454/merge_stmt_1532_PhiAck/$exit
      -- CP-element group 330: 	 branch_block_stmt_454/merge_stmt_1532_PhiAck/phi_stmt_1533_ack
      -- 
    phi_stmt_1533_ack_3777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1533_ack_0, ack => convolution3D_CP_1129_elements(330)); -- 
    req_2979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(330), ack => array_obj_ref_1565_index_offset_req_0); -- 
    req_2984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(330), ack => array_obj_ref_1565_index_offset_req_1); -- 
    req_2999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(330), ack => addr_of_1566_final_reg_req_1); -- 
    cr_3049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(330), ack => ptr_deref_1569_store_0_req_1); -- 
    -- CP-element group 331:  merge  fork  transition  place  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	213 
    -- CP-element group 331: 	232 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	233 
    -- CP-element group 331: 	234 
    -- CP-element group 331:  members (13) 
      -- CP-element group 331: 	 branch_block_stmt_454/merge_stmt_1573_PhiReqMerge
      -- CP-element group 331: 	 branch_block_stmt_454/merge_stmt_1573__exit__
      -- CP-element group 331: 	 branch_block_stmt_454/call_stmt_1576__entry__
      -- CP-element group 331: 	 branch_block_stmt_454/call_stmt_1576/$entry
      -- CP-element group 331: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_sample_start_
      -- CP-element group 331: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_update_start_
      -- CP-element group 331: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_Sample/$entry
      -- CP-element group 331: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_Sample/crr
      -- CP-element group 331: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_454/call_stmt_1576/call_stmt_1576_Update/ccr
      -- CP-element group 331: 	 branch_block_stmt_454/merge_stmt_1573_PhiAck/$entry
      -- CP-element group 331: 	 branch_block_stmt_454/merge_stmt_1573_PhiAck/$exit
      -- CP-element group 331: 	 branch_block_stmt_454/merge_stmt_1573_PhiAck/dummy
      -- 
    crr_3061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(331), ack => call_stmt_1576_call_req_0); -- 
    ccr_3066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(331), ack => call_stmt_1576_call_req_1); -- 
    convolution3D_CP_1129_elements(331) <= OrReduce(convolution3D_CP_1129_elements(213) & convolution3D_CP_1129_elements(232));
    -- CP-element group 332:  transition  output  delay-element  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	245 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	336 
    -- CP-element group 332:  members (5) 
      -- CP-element group 332: 	 branch_block_stmt_454/ifx_xend227_whilex_xbody_PhiReq/$exit
      -- CP-element group 332: 	 branch_block_stmt_454/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1644/$exit
      -- CP-element group 332: 	 branch_block_stmt_454/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/$exit
      -- CP-element group 332: 	 branch_block_stmt_454/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1650_konst_delay_trans
      -- CP-element group 332: 	 branch_block_stmt_454/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_req
      -- 
    phi_stmt_1644_req_3799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1644_req_3799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(332), ack => phi_stmt_1644_req_1); -- 
    -- Element group convolution3D_CP_1129_elements(332) is a control-delay.
    cp_element_332_delay: control_delay_element  generic map(name => " 332_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(245), ack => convolution3D_CP_1129_elements(332), clk => clk, reset =>reset);
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	261 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (2) 
      -- CP-element group 333: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/SplitProtocol/Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/SplitProtocol/Sample/ra
      -- 
    ra_3819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1647_inst_ack_0, ack => convolution3D_CP_1129_elements(333)); -- 
    -- CP-element group 334:  transition  input  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	261 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (2) 
      -- CP-element group 334: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/SplitProtocol/Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/SplitProtocol/Update/ca
      -- 
    ca_3824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1647_inst_ack_1, ack => convolution3D_CP_1129_elements(334)); -- 
    -- CP-element group 335:  join  transition  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 335: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/$exit
      -- CP-element group 335: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/$exit
      -- CP-element group 335: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/$exit
      -- CP-element group 335: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_sources/type_cast_1647/SplitProtocol/$exit
      -- CP-element group 335: 	 branch_block_stmt_454/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1644/phi_stmt_1644_req
      -- 
    phi_stmt_1644_req_3825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1644_req_3825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(335), ack => phi_stmt_1644_req_0); -- 
    convolution3D_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(333) & convolution3D_CP_1129_elements(334);
      gj_convolution3D_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  merge  transition  place  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	332 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (2) 
      -- CP-element group 336: 	 branch_block_stmt_454/merge_stmt_1643_PhiReqMerge
      -- CP-element group 336: 	 branch_block_stmt_454/merge_stmt_1643_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(336) <= OrReduce(convolution3D_CP_1129_elements(332) & convolution3D_CP_1129_elements(335));
    -- CP-element group 337:  fork  transition  place  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	246 
    -- CP-element group 337: 	247 
    -- CP-element group 337: 	248 
    -- CP-element group 337: 	250 
    -- CP-element group 337: 	251 
    -- CP-element group 337: 	252 
    -- CP-element group 337: 	253 
    -- CP-element group 337: 	256 
    -- CP-element group 337: 	257 
    -- CP-element group 337: 	258 
    -- CP-element group 337:  members (35) 
      -- CP-element group 337: 	 branch_block_stmt_454/merge_stmt_1643__exit__
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704__entry__
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_update_start_
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_Sample/rr
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1664_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/WPIPE_num_out_pipe_1666_Sample/req
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_update_start_
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_Sample/rr
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1671_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_update_start_
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_Sample/rr
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/type_cast_1675_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_update_start_
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1686_Update/ccr
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_update_start_
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_Sample/crr
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_454/assign_stmt_1656_to_assign_stmt_1704/call_stmt_1693_Update/ccr
      -- CP-element group 337: 	 branch_block_stmt_454/merge_stmt_1643_PhiAck/$exit
      -- CP-element group 337: 	 branch_block_stmt_454/merge_stmt_1643_PhiAck/phi_stmt_1644_ack
      -- 
    phi_stmt_1644_ack_3830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1644_ack_0, ack => convolution3D_CP_1129_elements(337)); -- 
    rr_3151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1664_inst_req_0); -- 
    cr_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1664_inst_req_1); -- 
    req_3165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => WPIPE_num_out_pipe_1666_inst_req_0); -- 
    rr_3179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1671_inst_req_0); -- 
    cr_3184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1671_inst_req_1); -- 
    rr_3193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1675_inst_req_0); -- 
    cr_3198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1675_inst_req_1); -- 
    ccr_3212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => call_stmt_1686_call_req_1); -- 
    crr_3221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => call_stmt_1693_call_req_0); -- 
    ccr_3226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => call_stmt_1693_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1144_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1422_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_953_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_1070 : std_logic_vector(63 downto 0);
    signal R_indvar355_1244_resized : std_logic_vector(13 downto 0);
    signal R_indvar355_1244_scaled : std_logic_vector(13 downto 0);
    signal R_indvar369_775_resized : std_logic_vector(13 downto 0);
    signal R_indvar369_775_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1091_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1091_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1564_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1564_scaled : std_logic_vector(13 downto 0);
    signal add102_821 : std_logic_vector(63 downto 0);
    signal add108_839 : std_logic_vector(63 downto 0);
    signal add114_857 : std_logic_vector(63 downto 0);
    signal add120_875 : std_logic_vector(63 downto 0);
    signal add1216x_xi312_1549 : std_logic_vector(63 downto 0);
    signal add1216x_xi_1076 : std_logic_vector(63 downto 0);
    signal add126_893 : std_logic_vector(63 downto 0);
    signal add132_911 : std_logic_vector(63 downto 0);
    signal add13_505 : std_logic_vector(15 downto 0);
    signal add171_1272 : std_logic_vector(63 downto 0);
    signal add177_1290 : std_logic_vector(63 downto 0);
    signal add183_1308 : std_logic_vector(63 downto 0);
    signal add189_1326 : std_logic_vector(63 downto 0);
    signal add195_1344 : std_logic_vector(63 downto 0);
    signal add201_1362 : std_logic_vector(63 downto 0);
    signal add207_1380 : std_logic_vector(63 downto 0);
    signal add23_530 : std_logic_vector(15 downto 0);
    signal add33_555 : std_logic_vector(15 downto 0);
    signal add43_580 : std_logic_vector(15 downto 0);
    signal add53_605 : std_logic_vector(15 downto 0);
    signal add63_630 : std_logic_vector(15 downto 0);
    signal add73_655 : std_logic_vector(15 downto 0);
    signal add96_803 : std_logic_vector(63 downto 0);
    signal add_480 : std_logic_vector(31 downto 0);
    signal addx_xi303_1510 : std_logic_vector(63 downto 0);
    signal addx_xi_1037 : std_logic_vector(63 downto 0);
    signal and217_1440 : std_logic_vector(63 downto 0);
    signal and264_1682 : std_logic_vector(7 downto 0);
    signal and_971 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1092_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1092_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1092_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1092_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1092_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1092_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1245_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1245_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1245_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1245_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1245_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1245_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1565_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1565_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1565_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1565_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1565_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1565_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_776_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_776_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_776_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_776_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_776_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_776_root_address : std_logic_vector(13 downto 0);
    signal arrayidx143_1094 : std_logic_vector(31 downto 0);
    signal arrayidx211_1247 : std_logic_vector(31 downto 0);
    signal arrayidx226_1567 : std_logic_vector(31 downto 0);
    signal arrayidx_778 : std_logic_vector(31 downto 0);
    signal call105_830 : std_logic_vector(7 downto 0);
    signal call111_848 : std_logic_vector(7 downto 0);
    signal call117_866 : std_logic_vector(7 downto 0);
    signal call11_496 : std_logic_vector(7 downto 0);
    signal call123_884 : std_logic_vector(7 downto 0);
    signal call129_902 : std_logic_vector(7 downto 0);
    signal call164_1250 : std_logic_vector(7 downto 0);
    signal call168_1263 : std_logic_vector(7 downto 0);
    signal call16_508 : std_logic_vector(7 downto 0);
    signal call174_1281 : std_logic_vector(7 downto 0);
    signal call180_1299 : std_logic_vector(7 downto 0);
    signal call186_1317 : std_logic_vector(7 downto 0);
    signal call192_1335 : std_logic_vector(7 downto 0);
    signal call198_1353 : std_logic_vector(7 downto 0);
    signal call204_1371 : std_logic_vector(7 downto 0);
    signal call21_521 : std_logic_vector(7 downto 0);
    signal call229_1576 : std_logic_vector(63 downto 0);
    signal call26_533 : std_logic_vector(7 downto 0);
    signal call288_1719 : std_logic_vector(63 downto 0);
    signal call2_471 : std_logic_vector(7 downto 0);
    signal call31_546 : std_logic_vector(7 downto 0);
    signal call36_558 : std_logic_vector(7 downto 0);
    signal call41_571 : std_logic_vector(7 downto 0);
    signal call46_583 : std_logic_vector(7 downto 0);
    signal call51_596 : std_logic_vector(7 downto 0);
    signal call56_608 : std_logic_vector(7 downto 0);
    signal call61_621 : std_logic_vector(7 downto 0);
    signal call66_633 : std_logic_vector(7 downto 0);
    signal call6_483 : std_logic_vector(7 downto 0);
    signal call71_646 : std_logic_vector(7 downto 0);
    signal call89_781 : std_logic_vector(7 downto 0);
    signal call93_794 : std_logic_vector(7 downto 0);
    signal call99_812 : std_logic_vector(7 downto 0);
    signal call_458 : std_logic_vector(7 downto 0);
    signal callx_xi301_1501 : std_logic_vector(7 downto 0);
    signal callx_xi_1028 : std_logic_vector(7 downto 0);
    signal cmp161321_1152 : std_logic_vector(0 downto 0);
    signal cmp325_685 : std_logic_vector(0 downto 0);
    signal cmpx_xi306_1525 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1052 : std_logic_vector(0 downto 0);
    signal conv101_816 : std_logic_vector(63 downto 0);
    signal conv107_834 : std_logic_vector(63 downto 0);
    signal conv113_852 : std_logic_vector(63 downto 0);
    signal conv119_870 : std_logic_vector(63 downto 0);
    signal conv125_888 : std_logic_vector(63 downto 0);
    signal conv12_500 : std_logic_vector(15 downto 0);
    signal conv131_906 : std_logic_vector(63 downto 0);
    signal conv145_1104 : std_logic_vector(63 downto 0);
    signal conv147_1108 : std_logic_vector(63 downto 0);
    signal conv150_1112 : std_logic_vector(63 downto 0);
    signal conv153_1116 : std_logic_vector(63 downto 0);
    signal conv155_1146 : std_logic_vector(63 downto 0);
    signal conv165_1254 : std_logic_vector(63 downto 0);
    signal conv170_1267 : std_logic_vector(63 downto 0);
    signal conv176_1285 : std_logic_vector(63 downto 0);
    signal conv182_1303 : std_logic_vector(63 downto 0);
    signal conv188_1321 : std_logic_vector(63 downto 0);
    signal conv194_1339 : std_logic_vector(63 downto 0);
    signal conv19_512 : std_logic_vector(15 downto 0);
    signal conv1_462 : std_logic_vector(31 downto 0);
    signal conv200_1357 : std_logic_vector(63 downto 0);
    signal conv206_1375 : std_logic_vector(63 downto 0);
    signal conv22_525 : std_logic_vector(15 downto 0);
    signal conv230_1716 : std_logic_vector(63 downto 0);
    signal conv255_1672 : std_logic_vector(63 downto 0);
    signal conv261_1676 : std_logic_vector(63 downto 0);
    signal conv263_1665 : std_logic_vector(7 downto 0);
    signal conv289_1724 : std_logic_vector(63 downto 0);
    signal conv29_537 : std_logic_vector(15 downto 0);
    signal conv2x_xi296_1463 : std_logic_vector(31 downto 0);
    signal conv2x_xi_990 : std_logic_vector(31 downto 0);
    signal conv32_550 : std_logic_vector(15 downto 0);
    signal conv39_562 : std_logic_vector(15 downto 0);
    signal conv3_475 : std_logic_vector(31 downto 0);
    signal conv42_575 : std_logic_vector(15 downto 0);
    signal conv49_587 : std_logic_vector(15 downto 0);
    signal conv52_600 : std_logic_vector(15 downto 0);
    signal conv59_612 : std_logic_vector(15 downto 0);
    signal conv5x_xi302_1505 : std_logic_vector(63 downto 0);
    signal conv5x_xi_1032 : std_logic_vector(63 downto 0);
    signal conv62_625 : std_logic_vector(15 downto 0);
    signal conv69_637 : std_logic_vector(15 downto 0);
    signal conv72_650 : std_logic_vector(15 downto 0);
    signal conv79_659 : std_logic_vector(31 downto 0);
    signal conv81_663 : std_logic_vector(31 downto 0);
    signal conv83_679 : std_logic_vector(63 downto 0);
    signal conv90_785 : std_logic_vector(63 downto 0);
    signal conv95_798 : std_logic_vector(63 downto 0);
    signal conv9_487 : std_logic_vector(15 downto 0);
    signal convx_xi305_1520 : std_logic_vector(31 downto 0);
    signal convx_xi_1047 : std_logic_vector(31 downto 0);
    signal elementx_x021x_xi300_1479 : std_logic_vector(63 downto 0);
    signal elementx_x021x_xi_1006 : std_logic_vector(63 downto 0);
    signal exitcond33_926 : std_logic_vector(0 downto 0);
    signal exitcond5_1704 : std_logic_vector(0 downto 0);
    signal exitcond_1395 : std_logic_vector(0 downto 0);
    signal iNsTr_35_1025 : std_logic_vector(15 downto 0);
    signal iNsTr_55_1459 : std_logic_vector(63 downto 0);
    signal iNsTr_65_1498 : std_logic_vector(15 downto 0);
    signal iNsTr_73_1543 : std_logic_vector(63 downto 0);
    signal indvar355_1233 : std_logic_vector(63 downto 0);
    signal indvar369_764 : std_logic_vector(63 downto 0);
    signal indvar_1644 : std_logic_vector(31 downto 0);
    signal indvarx_xnext356_1390 : std_logic_vector(63 downto 0);
    signal indvarx_xnext370_921 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1699 : std_logic_vector(31 downto 0);
    signal ix_x0x_xlcssa_958 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_1427 : std_logic_vector(63 downto 0);
    signal mul148_1121 : std_logic_vector(63 downto 0);
    signal mul151_1126 : std_logic_vector(63 downto 0);
    signal mul154_1131 : std_logic_vector(63 downto 0);
    signal mul236_1582 : std_logic_vector(15 downto 0);
    signal mul249_1595 : std_logic_vector(15 downto 0);
    signal mul254_1656 : std_logic_vector(31 downto 0);
    signal mul260_1661 : std_logic_vector(31 downto 0);
    signal mul82_673 : std_logic_vector(31 downto 0);
    signal mul_668 : std_logic_vector(31 downto 0);
    signal nx_x022x_xi299_1472 : std_logic_vector(15 downto 0);
    signal nx_x022x_xi_999 : std_logic_vector(15 downto 0);
    signal phitmp329_1424 : std_logic_vector(63 downto 0);
    signal phitmp_955 : std_logic_vector(63 downto 0);
    signal ptr_deref_1096_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1096_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1096_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1096_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1096_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1096_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1382_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1382_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1382_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1382_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1382_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1382_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1569_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1569_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1569_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1569_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1569_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1569_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_913_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_913_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_913_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_913_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_913_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_913_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext_1137 : std_logic_vector(63 downto 0);
    signal sh_promx_xi313_1555 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1082 : std_logic_vector(63 downto 0);
    signal shl104_827 : std_logic_vector(63 downto 0);
    signal shl10_493 : std_logic_vector(15 downto 0);
    signal shl110_845 : std_logic_vector(63 downto 0);
    signal shl116_863 : std_logic_vector(63 downto 0);
    signal shl122_881 : std_logic_vector(63 downto 0);
    signal shl128_899 : std_logic_vector(63 downto 0);
    signal shl14x_xi314_1560 : std_logic_vector(63 downto 0);
    signal shl14x_xi_1087 : std_logic_vector(63 downto 0);
    signal shl167_1260 : std_logic_vector(63 downto 0);
    signal shl173_1278 : std_logic_vector(63 downto 0);
    signal shl179_1296 : std_logic_vector(63 downto 0);
    signal shl185_1314 : std_logic_vector(63 downto 0);
    signal shl191_1332 : std_logic_vector(63 downto 0);
    signal shl197_1350 : std_logic_vector(63 downto 0);
    signal shl203_1368 : std_logic_vector(63 downto 0);
    signal shl20_518 : std_logic_vector(15 downto 0);
    signal shl30_543 : std_logic_vector(15 downto 0);
    signal shl40_568 : std_logic_vector(15 downto 0);
    signal shl50_593 : std_logic_vector(15 downto 0);
    signal shl60_618 : std_logic_vector(15 downto 0);
    signal shl70_643 : std_logic_vector(15 downto 0);
    signal shl8x_xi304_1516 : std_logic_vector(63 downto 0);
    signal shl8x_xi304x_xlcssa_1533 : std_logic_vector(63 downto 0);
    signal shl8x_xi_1043 : std_logic_vector(63 downto 0);
    signal shl8x_xix_xlcssa_1060 : std_logic_vector(63 downto 0);
    signal shl92_791 : std_logic_vector(63 downto 0);
    signal shl98_809 : std_logic_vector(63 downto 0);
    signal shl_468 : std_logic_vector(31 downto 0);
    signal shlx_xi297_1469 : std_logic_vector(31 downto 0);
    signal shlx_xi_996 : std_logic_vector(31 downto 0);
    signal sub273_1607 : std_logic_vector(15 downto 0);
    signal sub293_1729 : std_logic_vector(63 downto 0);
    signal sub_1601 : std_logic_vector(15 downto 0);
    signal tmp13_1175 : std_logic_vector(63 downto 0);
    signal tmp14_1179 : std_logic_vector(63 downto 0);
    signal tmp15_1184 : std_logic_vector(63 downto 0);
    signal tmp16_1188 : std_logic_vector(63 downto 0);
    signal tmp17_1193 : std_logic_vector(63 downto 0);
    signal tmp18_1197 : std_logic_vector(63 downto 0);
    signal tmp19_1202 : std_logic_vector(63 downto 0);
    signal tmp20_1206 : std_logic_vector(31 downto 0);
    signal tmp21_1211 : std_logic_vector(63 downto 0);
    signal tmp22_1217 : std_logic_vector(63 downto 0);
    signal tmp23_1223 : std_logic_vector(0 downto 0);
    signal tmp25_723 : std_logic_vector(31 downto 0);
    signal tmp26_728 : std_logic_vector(31 downto 0);
    signal tmp27_732 : std_logic_vector(31 downto 0);
    signal tmp28_737 : std_logic_vector(31 downto 0);
    signal tmp29_742 : std_logic_vector(63 downto 0);
    signal tmp30_748 : std_logic_vector(63 downto 0);
    signal tmp31_754 : std_logic_vector(0 downto 0);
    signal tmp330_1492 : std_logic_vector(15 downto 0);
    signal tmp331_1613 : std_logic_vector(15 downto 0);
    signal tmp350_1165 : std_logic_vector(63 downto 0);
    signal tmp351_1171 : std_logic_vector(0 downto 0);
    signal tmp352_1415 : std_logic_vector(63 downto 0);
    signal tmp359_697 : std_logic_vector(31 downto 0);
    signal tmp361_702 : std_logic_vector(31 downto 0);
    signal tmp362_707 : std_logic_vector(63 downto 0);
    signal tmp363_713 : std_logic_vector(63 downto 0);
    signal tmp364_719 : std_logic_vector(0 downto 0);
    signal tmp366_946 : std_logic_vector(63 downto 0);
    signal tmp3_1617 : std_logic_vector(31 downto 0);
    signal tmp4_1623 : std_logic_vector(31 downto 0);
    signal tmp6_1627 : std_logic_vector(31 downto 0);
    signal tmp7_1632 : std_logic_vector(15 downto 0);
    signal tmp8_1636 : std_logic_vector(31 downto 0);
    signal tmp9_1641 : std_logic_vector(31 downto 0);
    signal tmp_1019 : std_logic_vector(15 downto 0);
    signal tobool218_1446 : std_logic_vector(0 downto 0);
    signal tobool_977 : std_logic_vector(0 downto 0);
    signal type_cast_1003_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1005_wire : std_logic_vector(15 downto 0);
    signal type_cast_1010_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1012_wire : std_logic_vector(63 downto 0);
    signal type_cast_1017_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1023_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1041_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1063_wire : std_logic_vector(63 downto 0);
    signal type_cast_1068_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1074_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1080_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1135_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1140_wire : std_logic_vector(63 downto 0);
    signal type_cast_1143_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1150_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1163_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1169_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1209_wire : std_logic_vector(63 downto 0);
    signal type_cast_1215_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1221_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1228_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1237_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1239_wire : std_logic_vector(63 downto 0);
    signal type_cast_1258_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1276_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1294_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1312_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1330_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1348_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1366_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1388_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1407_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1413_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1418_wire : std_logic_vector(63 downto 0);
    signal type_cast_1421_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1430_wire : std_logic_vector(63 downto 0);
    signal type_cast_1433_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1438_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1444_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1467_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1476_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1478_wire : std_logic_vector(15 downto 0);
    signal type_cast_1483_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1485_wire : std_logic_vector(63 downto 0);
    signal type_cast_1490_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1496_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1514_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1536_wire : std_logic_vector(63 downto 0);
    signal type_cast_1541_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1547_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1553_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1585_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1589_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1599_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1605_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1611_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1621_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1647_wire : std_logic_vector(31 downto 0);
    signal type_cast_1650_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1680_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1697_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1714_wire : std_logic_vector(63 downto 0);
    signal type_cast_1722_wire : std_logic_vector(63 downto 0);
    signal type_cast_466_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_491_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_516_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_541_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_591_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_616_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_641_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_677_wire : std_logic_vector(63 downto 0);
    signal type_cast_683_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_705_wire : std_logic_vector(63 downto 0);
    signal type_cast_711_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_717_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_740_wire : std_logic_vector(63 downto 0);
    signal type_cast_746_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_752_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_759_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_767_wire : std_logic_vector(63 downto 0);
    signal type_cast_770_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_789_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_807_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_825_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_843_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_861_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_879_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_897_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_919_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_938_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_944_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_949_wire : std_logic_vector(63 downto 0);
    signal type_cast_952_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_961_wire : std_logic_vector(63 downto 0);
    signal type_cast_964_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_969_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_975_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_988_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_994_wire_constant : std_logic_vector(31 downto 0);
    signal umax24_1230 : std_logic_vector(63 downto 0);
    signal umax32_761 : std_logic_vector(63 downto 0);
    signal umax365_940 : std_logic_vector(63 downto 0);
    signal umax_1409 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1092_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1092_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1092_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1092_resized_base_address <= "00000000000000";
    array_obj_ref_1245_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1245_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1245_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1245_resized_base_address <= "00000000000000";
    array_obj_ref_1565_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1565_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1565_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1565_resized_base_address <= "00000000000000";
    array_obj_ref_776_constant_part_of_offset <= "00000000000000";
    array_obj_ref_776_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_776_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_776_resized_base_address <= "00000000000000";
    ptr_deref_1096_word_offset_0 <= "00000000000000";
    ptr_deref_1382_word_offset_0 <= "00000000000000";
    ptr_deref_1569_word_offset_0 <= "00000000000000";
    ptr_deref_913_word_offset_0 <= "00000000000000";
    type_cast_1003_wire_constant <= "0000000000000000";
    type_cast_1010_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1017_wire_constant <= "0000000000000001";
    type_cast_1023_wire_constant <= "0000000000000001";
    type_cast_1041_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1068_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1074_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1080_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1135_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1143_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1150_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1163_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1169_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1215_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1221_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1228_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1237_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1258_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1276_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1294_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1312_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1330_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1348_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1366_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1388_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1407_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1413_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1421_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1433_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1438_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1444_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1457_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1467_wire_constant <= "00000000000000000000000000000110";
    type_cast_1476_wire_constant <= "0000000000000000";
    type_cast_1483_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1490_wire_constant <= "0000000000000001";
    type_cast_1496_wire_constant <= "0000000000000001";
    type_cast_1514_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1541_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1547_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1553_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1585_wire_constant <= "11001000";
    type_cast_1589_wire_constant <= "11001000";
    type_cast_1599_wire_constant <= "1111111111111111";
    type_cast_1605_wire_constant <= "1111111111111111";
    type_cast_1611_wire_constant <= "1111111111111111";
    type_cast_1621_wire_constant <= "00000000000000000000000000000001";
    type_cast_1650_wire_constant <= "00000000000000000000000000000000";
    type_cast_1680_wire_constant <= "00000001";
    type_cast_1697_wire_constant <= "00000000000000000000000000000001";
    type_cast_466_wire_constant <= "00000000000000000000000000001000";
    type_cast_491_wire_constant <= "0000000000001000";
    type_cast_516_wire_constant <= "0000000000001000";
    type_cast_541_wire_constant <= "0000000000001000";
    type_cast_566_wire_constant <= "0000000000001000";
    type_cast_591_wire_constant <= "0000000000001000";
    type_cast_616_wire_constant <= "0000000000001000";
    type_cast_641_wire_constant <= "0000000000001000";
    type_cast_683_wire_constant <= "00000000000000000000000000000011";
    type_cast_711_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_717_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_746_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_752_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_759_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_770_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_789_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_807_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_825_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_843_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_861_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_879_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_897_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_919_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_938_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_944_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_952_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_964_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_969_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_975_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_988_wire_constant <= "00000000000000000000000000000001";
    type_cast_994_wire_constant <= "00000000000000000000000000000110";
    phi_stmt_1006: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1010_wire_constant & type_cast_1012_wire;
      req <= phi_stmt_1006_req_0 & phi_stmt_1006_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1006",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1006_ack_0,
          idata => idata,
          odata => elementx_x021x_xi_1006,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1006
    phi_stmt_1060: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1063_wire;
      req(0) <= phi_stmt_1060_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1060",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1060_ack_0,
          idata => idata,
          odata => shl8x_xix_xlcssa_1060,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1060
    phi_stmt_1233: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1237_wire_constant & type_cast_1239_wire;
      req <= phi_stmt_1233_req_0 & phi_stmt_1233_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1233",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1233_ack_0,
          idata => idata,
          odata => indvar355_1233,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1233
    phi_stmt_1427: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1430_wire & type_cast_1433_wire_constant;
      req <= phi_stmt_1427_req_0 & phi_stmt_1427_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1427",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1427_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_1427,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1427
    phi_stmt_1472: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1476_wire_constant & type_cast_1478_wire;
      req <= phi_stmt_1472_req_0 & phi_stmt_1472_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1472",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1472_ack_0,
          idata => idata,
          odata => nx_x022x_xi299_1472,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1472
    phi_stmt_1479: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1483_wire_constant & type_cast_1485_wire;
      req <= phi_stmt_1479_req_0 & phi_stmt_1479_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1479",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1479_ack_0,
          idata => idata,
          odata => elementx_x021x_xi300_1479,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1479
    phi_stmt_1533: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1536_wire;
      req(0) <= phi_stmt_1533_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1533",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1533_ack_0,
          idata => idata,
          odata => shl8x_xi304x_xlcssa_1533,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1533
    phi_stmt_1644: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1647_wire & type_cast_1650_wire_constant;
      req <= phi_stmt_1644_req_0 & phi_stmt_1644_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1644",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1644_ack_0,
          idata => idata,
          odata => indvar_1644,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1644
    phi_stmt_764: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_767_wire & type_cast_770_wire_constant;
      req <= phi_stmt_764_req_0 & phi_stmt_764_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_764",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_764_ack_0,
          idata => idata,
          odata => indvar369_764,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_764
    phi_stmt_958: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_961_wire & type_cast_964_wire_constant;
      req <= phi_stmt_958_req_0 & phi_stmt_958_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_958",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_958_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_958,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_958
    phi_stmt_999: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1003_wire_constant & type_cast_1005_wire;
      req <= phi_stmt_999_req_0 & phi_stmt_999_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_999",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_999_ack_0,
          idata => idata,
          odata => nx_x022x_xi_999,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_999
    -- flow-through select operator MUX_1229_inst
    umax24_1230 <= tmp22_1217 when (tmp23_1223(0) /=  '0') else type_cast_1228_wire_constant;
    -- flow-through select operator MUX_1408_inst
    umax_1409 <= tmp350_1165 when (tmp351_1171(0) /=  '0') else type_cast_1407_wire_constant;
    -- flow-through select operator MUX_760_inst
    umax32_761 <= tmp30_748 when (tmp31_754(0) /=  '0') else type_cast_759_wire_constant;
    -- flow-through select operator MUX_939_inst
    umax365_940 <= tmp363_713 when (tmp364_719(0) /=  '0') else type_cast_938_wire_constant;
    addr_of_1093_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1093_final_reg_req_0;
      addr_of_1093_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1093_final_reg_req_1;
      addr_of_1093_final_reg_ack_1<= rack(0);
      addr_of_1093_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1093_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1092_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx143_1094,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1246_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1246_final_reg_req_0;
      addr_of_1246_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1246_final_reg_req_1;
      addr_of_1246_final_reg_ack_1<= rack(0);
      addr_of_1246_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1246_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1245_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx211_1247,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1566_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1566_final_reg_req_0;
      addr_of_1566_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1566_final_reg_req_1;
      addr_of_1566_final_reg_ack_1<= rack(0);
      addr_of_1566_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1566_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1565_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx226_1567,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_777_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_777_final_reg_req_0;
      addr_of_777_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_777_final_reg_req_1;
      addr_of_777_final_reg_ack_1<= rack(0);
      addr_of_777_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_777_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_776_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_778,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1005_inst_req_0;
      type_cast_1005_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1005_inst_req_1;
      type_cast_1005_inst_ack_1<= rack(0);
      type_cast_1005_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1005_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_35_1025,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1005_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1012_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1012_inst_req_0;
      type_cast_1012_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1012_inst_req_1;
      type_cast_1012_inst_ack_1<= rack(0);
      type_cast_1012_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1012_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1043,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1012_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1031_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1031_inst_req_0;
      type_cast_1031_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1031_inst_req_1;
      type_cast_1031_inst_ack_1<= rack(0);
      type_cast_1031_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1031_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1028,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_1032,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1046_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1046_inst_req_0;
      type_cast_1046_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1046_inst_req_1;
      type_cast_1046_inst_ack_1<= rack(0);
      type_cast_1046_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1046_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1019,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1047,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1063_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1063_inst_req_0;
      type_cast_1063_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1063_inst_req_1;
      type_cast_1063_inst_ack_1<= rack(0);
      type_cast_1063_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1063_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1043,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1063_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1103_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1103_inst_req_0;
      type_cast_1103_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1103_inst_req_1;
      type_cast_1103_inst_ack_1<= rack(0);
      type_cast_1103_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1103_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_530,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1104,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1107_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1107_inst_req_0;
      type_cast_1107_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1107_inst_req_1;
      type_cast_1107_inst_ack_1<= rack(0);
      type_cast_1107_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1107_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_655,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_1108,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1111_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1111_inst_req_0;
      type_cast_1111_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1111_inst_req_1;
      type_cast_1111_inst_ack_1<= rack(0);
      type_cast_1111_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1111_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv150_1112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1115_inst_req_0;
      type_cast_1115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1115_inst_req_1;
      type_cast_1115_inst_ack_1<= rack(0);
      type_cast_1115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1115_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1116,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1140_inst
    process(sext_1137) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1137(63 downto 0);
      type_cast_1140_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1145_inst
    process(ASHR_i64_i64_1144_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1144_wire(63 downto 0);
      conv155_1146 <= tmp_var; -- 
    end process;
    type_cast_1174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1174_inst_req_0;
      type_cast_1174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1174_inst_req_1;
      type_cast_1174_inst_ack_1<= rack(0);
      type_cast_1174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_1175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1178_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1178_inst_req_0;
      type_cast_1178_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1178_inst_req_1;
      type_cast_1178_inst_ack_1<= rack(0);
      type_cast_1178_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1178_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_530,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp14_1179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1187_inst_req_0;
      type_cast_1187_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1187_inst_req_1;
      type_cast_1187_inst_ack_1<= rack(0);
      type_cast_1187_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp16_1188,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1196_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1196_inst_req_0;
      type_cast_1196_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1196_inst_req_1;
      type_cast_1196_inst_ack_1<= rack(0);
      type_cast_1196_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1196_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_655,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp18_1197,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1205_inst_req_0;
      type_cast_1205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1205_inst_req_1;
      type_cast_1205_inst_ack_1<= rack(0);
      type_cast_1205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp19_1202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1210_inst_req_0;
      type_cast_1210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1210_inst_req_1;
      type_cast_1210_inst_ack_1<= rack(0);
      type_cast_1210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1209_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp21_1211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1239_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1239_inst_req_0;
      type_cast_1239_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1239_inst_req_1;
      type_cast_1239_inst_ack_1<= rack(0);
      type_cast_1239_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1239_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext356_1390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1239_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1253_inst_req_0;
      type_cast_1253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1253_inst_req_1;
      type_cast_1253_inst_ack_1<= rack(0);
      type_cast_1253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_1250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_1254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1266_inst_req_0;
      type_cast_1266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1266_inst_req_1;
      type_cast_1266_inst_ack_1<= rack(0);
      type_cast_1266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_1263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1284_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1284_inst_req_0;
      type_cast_1284_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1284_inst_req_1;
      type_cast_1284_inst_ack_1<= rack(0);
      type_cast_1284_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1284_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_1281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_1285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1302_inst_req_0;
      type_cast_1302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1302_inst_req_1;
      type_cast_1302_inst_ack_1<= rack(0);
      type_cast_1302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_1299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_1303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1320_inst_req_0;
      type_cast_1320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1320_inst_req_1;
      type_cast_1320_inst_ack_1<= rack(0);
      type_cast_1320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_1317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_1321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1338_inst_req_0;
      type_cast_1338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1338_inst_req_1;
      type_cast_1338_inst_ack_1<= rack(0);
      type_cast_1338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call192_1335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv194_1339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1356_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1356_inst_req_0;
      type_cast_1356_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1356_inst_req_1;
      type_cast_1356_inst_ack_1<= rack(0);
      type_cast_1356_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1356_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call198_1353,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_1357,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1374_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1374_inst_req_0;
      type_cast_1374_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1374_inst_req_1;
      type_cast_1374_inst_ack_1<= rack(0);
      type_cast_1374_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1374_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call204_1371,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_1375,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1418_inst
    process(tmp352_1415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp352_1415(63 downto 0);
      type_cast_1418_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1423_inst
    process(ASHR_i64_i64_1422_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1422_wire(63 downto 0);
      phitmp329_1424 <= tmp_var; -- 
    end process;
    type_cast_1430_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1430_inst_req_0;
      type_cast_1430_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1430_inst_req_1;
      type_cast_1430_inst_ack_1<= rack(0);
      type_cast_1430_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1430_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp329_1424,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1430_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1462_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1462_inst_req_0;
      type_cast_1462_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1462_inst_req_1;
      type_cast_1462_inst_ack_1<= rack(0);
      type_cast_1462_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1462_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_55_1459,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi296_1463,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1478_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1478_inst_req_0;
      type_cast_1478_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1478_inst_req_1;
      type_cast_1478_inst_ack_1<= rack(0);
      type_cast_1478_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1478_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_65_1498,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1478_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1485_inst_req_0;
      type_cast_1485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1485_inst_req_1;
      type_cast_1485_inst_ack_1<= rack(0);
      type_cast_1485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi304_1516,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1485_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1504_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1504_inst_req_0;
      type_cast_1504_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1504_inst_req_1;
      type_cast_1504_inst_ack_1<= rack(0);
      type_cast_1504_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1504_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi301_1501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi302_1505,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1519_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1519_inst_req_0;
      type_cast_1519_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1519_inst_req_1;
      type_cast_1519_inst_ack_1<= rack(0);
      type_cast_1519_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1519_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp330_1492,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi305_1520,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1536_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1536_inst_req_0;
      type_cast_1536_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1536_inst_req_1;
      type_cast_1536_inst_ack_1<= rack(0);
      type_cast_1536_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1536_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi304_1516,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1536_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1616_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1616_inst_req_0;
      type_cast_1616_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1616_inst_req_1;
      type_cast_1616_inst_ack_1<= rack(0);
      type_cast_1616_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1616_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp331_1613,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1617,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1626_inst_req_0;
      type_cast_1626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1626_inst_req_1;
      type_cast_1626_inst_ack_1<= rack(0);
      type_cast_1626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_1627,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1635_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1635_inst_req_0;
      type_cast_1635_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1635_inst_req_1;
      type_cast_1635_inst_ack_1<= rack(0);
      type_cast_1635_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1635_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp7_1632,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp8_1636,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1647_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1647_inst_req_0;
      type_cast_1647_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1647_inst_req_1;
      type_cast_1647_inst_ack_1<= rack(0);
      type_cast_1647_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1647_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1699,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1647_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1664_inst_req_0;
      type_cast_1664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1664_inst_req_1;
      type_cast_1664_inst_ack_1<= rack(0);
      type_cast_1664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvar_1644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv263_1665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1671_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1671_inst_req_0;
      type_cast_1671_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1671_inst_req_1;
      type_cast_1671_inst_ack_1<= rack(0);
      type_cast_1671_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1671_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul254_1656,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_1672,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1675_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1675_inst_req_0;
      type_cast_1675_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1675_inst_req_1;
      type_cast_1675_inst_ack_1<= rack(0);
      type_cast_1675_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1675_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul260_1661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv261_1676,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1715_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1715_inst_req_0;
      type_cast_1715_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1715_inst_req_1;
      type_cast_1715_inst_ack_1<= rack(0);
      type_cast_1715_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1715_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1714_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv230_1716,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1723_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1723_inst_req_0;
      type_cast_1723_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1723_inst_req_1;
      type_cast_1723_inst_ack_1<= rack(0);
      type_cast_1723_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1723_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1722_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv289_1724,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_461_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_461_inst_req_0;
      type_cast_461_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_461_inst_req_1;
      type_cast_461_inst_ack_1<= rack(0);
      type_cast_461_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_461_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_458,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_462,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_474_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_474_inst_req_0;
      type_cast_474_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_474_inst_req_1;
      type_cast_474_inst_ack_1<= rack(0);
      type_cast_474_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_474_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_471,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_475,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_486_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_486_inst_req_0;
      type_cast_486_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_486_inst_req_1;
      type_cast_486_inst_ack_1<= rack(0);
      type_cast_486_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_486_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_483,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_487,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_499_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_499_inst_req_0;
      type_cast_499_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_499_inst_req_1;
      type_cast_499_inst_ack_1<= rack(0);
      type_cast_499_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_499_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_496,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_500,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_511_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_511_inst_req_0;
      type_cast_511_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_511_inst_req_1;
      type_cast_511_inst_ack_1<= rack(0);
      type_cast_511_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_511_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_508,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_512,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_524_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_524_inst_req_0;
      type_cast_524_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_524_inst_req_1;
      type_cast_524_inst_ack_1<= rack(0);
      type_cast_524_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_524_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_521,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_525,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_536_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_536_inst_req_0;
      type_cast_536_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_536_inst_req_1;
      type_cast_536_inst_ack_1<= rack(0);
      type_cast_536_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_536_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_533,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_537,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_549_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_549_inst_req_0;
      type_cast_549_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_549_inst_req_1;
      type_cast_549_inst_ack_1<= rack(0);
      type_cast_549_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_549_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_546,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_550,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_561_inst_req_0;
      type_cast_561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_561_inst_req_1;
      type_cast_561_inst_ack_1<= rack(0);
      type_cast_561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_574_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_574_inst_req_0;
      type_cast_574_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_574_inst_req_1;
      type_cast_574_inst_ack_1<= rack(0);
      type_cast_574_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_574_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_571,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_575,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_586_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_586_inst_req_0;
      type_cast_586_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_586_inst_req_1;
      type_cast_586_inst_ack_1<= rack(0);
      type_cast_586_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_586_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_583,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_587,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_599_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_599_inst_req_0;
      type_cast_599_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_599_inst_req_1;
      type_cast_599_inst_ack_1<= rack(0);
      type_cast_599_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_599_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_596,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_600,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_611_inst_req_0;
      type_cast_611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_611_inst_req_1;
      type_cast_611_inst_ack_1<= rack(0);
      type_cast_611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_612,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_624_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_624_inst_req_0;
      type_cast_624_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_624_inst_req_1;
      type_cast_624_inst_ack_1<= rack(0);
      type_cast_624_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_624_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_621,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_625,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_636_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_636_inst_req_0;
      type_cast_636_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_636_inst_req_1;
      type_cast_636_inst_ack_1<= rack(0);
      type_cast_636_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_636_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_633,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_637,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_649_inst_req_0;
      type_cast_649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_649_inst_req_1;
      type_cast_649_inst_ack_1<= rack(0);
      type_cast_649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_658_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_658_inst_req_0;
      type_cast_658_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_658_inst_req_1;
      type_cast_658_inst_ack_1<= rack(0);
      type_cast_658_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_658_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_659,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_662_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_662_inst_req_0;
      type_cast_662_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_662_inst_req_1;
      type_cast_662_inst_ack_1<= rack(0);
      type_cast_662_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_662_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_530,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_663,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_678_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_678_inst_req_0;
      type_cast_678_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_678_inst_req_1;
      type_cast_678_inst_ack_1<= rack(0);
      type_cast_678_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_678_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_677_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_679,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_706_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_706_inst_req_0;
      type_cast_706_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_706_inst_req_1;
      type_cast_706_inst_ack_1<= rack(0);
      type_cast_706_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_706_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_705_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp362_707,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_722_inst_req_0;
      type_cast_722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_722_inst_req_1;
      type_cast_722_inst_ack_1<= rack(0);
      type_cast_722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp25_723,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_731_inst_req_0;
      type_cast_731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_731_inst_req_1;
      type_cast_731_inst_ack_1<= rack(0);
      type_cast_731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_530,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp27_732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_741_inst_req_0;
      type_cast_741_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_741_inst_req_1;
      type_cast_741_inst_ack_1<= rack(0);
      type_cast_741_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_741_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_740_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp29_742,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_767_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_767_inst_req_0;
      type_cast_767_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_767_inst_req_1;
      type_cast_767_inst_ack_1<= rack(0);
      type_cast_767_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_767_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext370_921,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_767_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_784_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_784_inst_req_0;
      type_cast_784_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_784_inst_req_1;
      type_cast_784_inst_ack_1<= rack(0);
      type_cast_784_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_784_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_781,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_785,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_797_inst_req_0;
      type_cast_797_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_797_inst_req_1;
      type_cast_797_inst_ack_1<= rack(0);
      type_cast_797_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_797_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_794,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_798,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_815_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_815_inst_req_0;
      type_cast_815_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_815_inst_req_1;
      type_cast_815_inst_ack_1<= rack(0);
      type_cast_815_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_815_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call99_812,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_816,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_833_inst_req_0;
      type_cast_833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_833_inst_req_1;
      type_cast_833_inst_ack_1<= rack(0);
      type_cast_833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call105_830,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_834,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_851_inst_req_0;
      type_cast_851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_851_inst_req_1;
      type_cast_851_inst_ack_1<= rack(0);
      type_cast_851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_848,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_869_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_869_inst_req_0;
      type_cast_869_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_869_inst_req_1;
      type_cast_869_inst_ack_1<= rack(0);
      type_cast_869_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_869_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call117_866,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_870,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_887_inst_req_0;
      type_cast_887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_887_inst_req_1;
      type_cast_887_inst_ack_1<= rack(0);
      type_cast_887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call123_884,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_905_inst_req_0;
      type_cast_905_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_905_inst_req_1;
      type_cast_905_inst_ack_1<= rack(0);
      type_cast_905_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_905_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_902,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_906,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_949_inst
    process(tmp366_946) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp366_946(63 downto 0);
      type_cast_949_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_954_inst
    process(ASHR_i64_i64_953_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_953_wire(63 downto 0);
      phitmp_955 <= tmp_var; -- 
    end process;
    type_cast_961_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_961_inst_req_0;
      type_cast_961_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_961_inst_req_1;
      type_cast_961_inst_ack_1<= rack(0);
      type_cast_961_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_961_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_955,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_961_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1092_index_1_rename
    process(R_ix_x0x_xlcssa_1091_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1091_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1091_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1092_index_1_resize
    process(ix_x0x_xlcssa_958) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_958;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1091_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1092_root_address_inst
    process(array_obj_ref_1092_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1092_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1092_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1245_index_1_rename
    process(R_indvar355_1244_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar355_1244_resized;
      ov(13 downto 0) := iv;
      R_indvar355_1244_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1245_index_1_resize
    process(indvar355_1233) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar355_1233;
      ov := iv(13 downto 0);
      R_indvar355_1244_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1245_root_address_inst
    process(array_obj_ref_1245_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1245_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1245_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1565_index_1_rename
    process(R_ix_x1x_xlcssa_1564_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_1564_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_1564_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1565_index_1_resize
    process(ix_x1x_xlcssa_1427) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_1427;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_1564_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1565_root_address_inst
    process(array_obj_ref_1565_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1565_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1565_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_776_index_1_rename
    process(R_indvar369_775_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar369_775_resized;
      ov(13 downto 0) := iv;
      R_indvar369_775_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_776_index_1_resize
    process(indvar369_764) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar369_764;
      ov := iv(13 downto 0);
      R_indvar369_775_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_776_root_address_inst
    process(array_obj_ref_776_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_776_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_776_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_addr_0
    process(ptr_deref_1096_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1096_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1096_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_base_resize
    process(arrayidx143_1094) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx143_1094;
      ov := iv(13 downto 0);
      ptr_deref_1096_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_gather_scatter
    process(shl14x_xi_1087) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi_1087;
      ov(63 downto 0) := iv;
      ptr_deref_1096_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_root_address_inst
    process(ptr_deref_1096_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1096_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1096_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1382_addr_0
    process(ptr_deref_1382_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1382_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1382_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1382_base_resize
    process(arrayidx211_1247) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx211_1247;
      ov := iv(13 downto 0);
      ptr_deref_1382_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1382_gather_scatter
    process(add207_1380) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add207_1380;
      ov(63 downto 0) := iv;
      ptr_deref_1382_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1382_root_address_inst
    process(ptr_deref_1382_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1382_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1382_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1569_addr_0
    process(ptr_deref_1569_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1569_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1569_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1569_base_resize
    process(arrayidx226_1567) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx226_1567;
      ov := iv(13 downto 0);
      ptr_deref_1569_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1569_gather_scatter
    process(shl14x_xi314_1560) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi314_1560;
      ov(63 downto 0) := iv;
      ptr_deref_1569_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1569_root_address_inst
    process(ptr_deref_1569_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1569_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1569_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_addr_0
    process(ptr_deref_913_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_913_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_913_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_base_resize
    process(arrayidx_778) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_778;
      ov := iv(13 downto 0);
      ptr_deref_913_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_gather_scatter
    process(add132_911) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add132_911;
      ov(63 downto 0) := iv;
      ptr_deref_913_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_root_address_inst
    process(ptr_deref_913_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_913_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_913_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1053_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_1052;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1053_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1053_branch_req_0,
          ack0 => if_stmt_1053_branch_ack_0,
          ack1 => if_stmt_1053_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1153_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp161321_1152;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1153_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1153_branch_req_0,
          ack0 => if_stmt_1153_branch_ack_0,
          ack1 => if_stmt_1153_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1396_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1395;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1396_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1396_branch_req_0,
          ack0 => if_stmt_1396_branch_ack_0,
          ack1 => if_stmt_1396_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1447_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool218_1446;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1447_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1447_branch_req_0,
          ack0 => if_stmt_1447_branch_ack_0,
          ack1 => if_stmt_1447_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1526_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi306_1525;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1526_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1526_branch_req_0,
          ack0 => if_stmt_1526_branch_ack_0,
          ack1 => if_stmt_1526_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1705_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_1704;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1705_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1705_branch_req_0,
          ack0 => if_stmt_1705_branch_ack_0,
          ack1 => if_stmt_1705_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_686_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp325_685;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_686_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_686_branch_req_0,
          ack0 => if_stmt_686_branch_ack_0,
          ack1 => if_stmt_686_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_927_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond33_926;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_927_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_927_branch_req_0,
          ack0 => if_stmt_927_branch_ack_0,
          ack1 => if_stmt_927_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_978_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_977;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_978_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_978_branch_req_0,
          ack0 => if_stmt_978_branch_ack_0,
          ack1 => if_stmt_978_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1018_inst
    process(nx_x022x_xi_999) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_999, type_cast_1017_wire_constant, tmp_var);
      tmp_1019 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1024_inst
    process(nx_x022x_xi_999) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_999, type_cast_1023_wire_constant, tmp_var);
      iNsTr_35_1025 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1491_inst
    process(nx_x022x_xi299_1472) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi299_1472, type_cast_1490_wire_constant, tmp_var);
      tmp330_1492 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1497_inst
    process(nx_x022x_xi299_1472) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi299_1472, type_cast_1496_wire_constant, tmp_var);
      iNsTr_65_1498 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1600_inst
    process(add43_580) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add43_580, type_cast_1599_wire_constant, tmp_var);
      sub_1601 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1606_inst
    process(add63_630) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add63_630, type_cast_1605_wire_constant, tmp_var);
      sub273_1607 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1612_inst
    process(add53_605) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_605, type_cast_1611_wire_constant, tmp_var);
      tmp331_1613 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1622_inst
    process(tmp3_1617) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1617, type_cast_1621_wire_constant, tmp_var);
      tmp4_1623 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1660_inst
    process(tmp9_1641, mul254_1656) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp9_1641, mul254_1656, tmp_var);
      mul260_1661 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1698_inst
    process(indvar_1644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1644, type_cast_1697_wire_constant, tmp_var);
      indvarx_xnext_1699 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1389_inst
    process(indvar355_1233) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar355_1233, type_cast_1388_wire_constant, tmp_var);
      indvarx_xnext356_1390 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_920_inst
    process(indvar369_764) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar369_764, type_cast_919_wire_constant, tmp_var);
      indvarx_xnext370_921 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1468_inst
    process(conv2x_xi296_1463) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi296_1463, type_cast_1467_wire_constant, tmp_var);
      shlx_xi297_1469 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_995_inst
    process(conv2x_xi_990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_990, type_cast_994_wire_constant, tmp_var);
      shlx_xi_996 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1075_inst
    process(Bx_xnot_1070) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_1070, type_cast_1074_wire_constant, tmp_var);
      add1216x_xi_1076 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1439_inst
    process(conv155_1146) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv155_1146, type_cast_1438_wire_constant, tmp_var);
      and217_1440 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1548_inst
    process(iNsTr_73_1543) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_73_1543, type_cast_1547_wire_constant, tmp_var);
      add1216x_xi312_1549 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_970_inst
    process(conv83_679) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv83_679, type_cast_969_wire_constant, tmp_var);
      and_971 <= tmp_var; --
    end process;
    -- binary operator AND_u8_u8_1681_inst
    process(conv263_1665) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv263_1665, type_cast_1680_wire_constant, tmp_var);
      and264_1682 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1144_inst
    process(type_cast_1140_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1140_wire, type_cast_1143_wire_constant, tmp_var);
      ASHR_i64_i64_1144_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1422_inst
    process(type_cast_1418_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1418_wire, type_cast_1421_wire_constant, tmp_var);
      ASHR_i64_i64_1422_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_953_inst
    process(type_cast_949_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_949_wire, type_cast_952_wire_constant, tmp_var);
      ASHR_i64_i64_953_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1703_inst
    process(indvarx_xnext_1699, tmp4_1623) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1699, tmp4_1623, tmp_var);
      exitcond5_1704 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1394_inst
    process(indvarx_xnext356_1390, umax24_1230) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext356_1390, umax24_1230, tmp_var);
      exitcond_1395 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1445_inst
    process(and217_1440) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and217_1440, type_cast_1444_wire_constant, tmp_var);
      tobool218_1446 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_925_inst
    process(indvarx_xnext370_921, umax32_761) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext370_921, umax32_761, tmp_var);
      exitcond33_926 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_976_inst
    process(and_971) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_971, type_cast_975_wire_constant, tmp_var);
      tobool_977 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1164_inst
    process(conv155_1146) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_1146, type_cast_1163_wire_constant, tmp_var);
      tmp350_1165 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1216_inst
    process(tmp21_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp21_1211, type_cast_1215_wire_constant, tmp_var);
      tmp22_1217 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_712_inst
    process(tmp362_707) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp362_707, type_cast_711_wire_constant, tmp_var);
      tmp363_713 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_747_inst
    process(tmp29_742) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp29_742, type_cast_746_wire_constant, tmp_var);
      tmp30_748 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1581_inst
    process(add73_655, add23_530) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_655, add23_530, tmp_var);
      mul236_1582 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1594_inst
    process(add43_580, add33_555) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add43_580, add33_555, tmp_var);
      mul249_1595 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1631_inst
    process(add73_655, add23_530) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_655, add23_530, tmp_var);
      tmp7_1632 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1640_inst
    process(tmp6_1627, tmp8_1636) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp6_1627, tmp8_1636, tmp_var);
      tmp9_1641 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1655_inst
    process(tmp9_1641, indvar_1644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp9_1641, indvar_1644, tmp_var);
      mul254_1656 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_667_inst
    process(conv79_659, add_480) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_659, add_480, tmp_var);
      mul_668 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_672_inst
    process(mul_668, conv81_663) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_668, conv81_663, tmp_var);
      mul82_673 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_696_inst
    process(add_480, conv79_659) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_480, conv79_659, tmp_var);
      tmp359_697 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_701_inst
    process(tmp359_697, conv81_663) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp359_697, conv81_663, tmp_var);
      tmp361_702 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_727_inst
    process(add_480, tmp25_723) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_480, tmp25_723, tmp_var);
      tmp26_728 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_736_inst
    process(tmp26_728, tmp27_732) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp26_728, tmp27_732, tmp_var);
      tmp28_737 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1120_inst
    process(conv153_1116, conv145_1104) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv153_1116, conv145_1104, tmp_var);
      mul148_1121 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1125_inst
    process(mul148_1121, conv150_1112) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul148_1121, conv150_1112, tmp_var);
      mul151_1126 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1130_inst
    process(mul151_1126, conv147_1108) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul151_1126, conv147_1108, tmp_var);
      mul154_1131 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1183_inst
    process(tmp13_1175, tmp14_1179) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_1175, tmp14_1179, tmp_var);
      tmp15_1184 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1192_inst
    process(tmp15_1184, tmp16_1188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp15_1184, tmp16_1188, tmp_var);
      tmp17_1193 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1201_inst
    process(tmp17_1193, tmp18_1197) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp17_1193, tmp18_1197, tmp_var);
      tmp19_1202 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_504_inst
    process(shl10_493, conv12_500) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_493, conv12_500, tmp_var);
      add13_505 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_529_inst
    process(shl20_518, conv22_525) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_518, conv22_525, tmp_var);
      add23_530 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_554_inst
    process(shl30_543, conv32_550) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_543, conv32_550, tmp_var);
      add33_555 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_579_inst
    process(shl40_568, conv42_575) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_568, conv42_575, tmp_var);
      add43_580 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_604_inst
    process(shl50_593, conv52_600) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_593, conv52_600, tmp_var);
      add53_605 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_629_inst
    process(shl60_618, conv62_625) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_618, conv62_625, tmp_var);
      add63_630 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_654_inst
    process(shl70_643, conv72_650) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_643, conv72_650, tmp_var);
      add73_655 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_479_inst
    process(shl_468, conv3_475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_468, conv3_475, tmp_var);
      add_480 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1036_inst
    process(conv5x_xi_1032, elementx_x021x_xi_1006) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_1032, elementx_x021x_xi_1006, tmp_var);
      addx_xi_1037 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1271_inst
    process(shl167_1260, conv170_1267) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_1260, conv170_1267, tmp_var);
      add171_1272 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1289_inst
    process(shl173_1278, conv176_1285) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_1278, conv176_1285, tmp_var);
      add177_1290 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1307_inst
    process(shl179_1296, conv182_1303) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl179_1296, conv182_1303, tmp_var);
      add183_1308 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1325_inst
    process(shl185_1314, conv188_1321) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl185_1314, conv188_1321, tmp_var);
      add189_1326 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1343_inst
    process(shl191_1332, conv194_1339) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl191_1332, conv194_1339, tmp_var);
      add195_1344 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1361_inst
    process(shl197_1350, conv200_1357) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl197_1350, conv200_1357, tmp_var);
      add201_1362 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1379_inst
    process(shl203_1368, conv206_1375) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl203_1368, conv206_1375, tmp_var);
      add207_1380 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1509_inst
    process(conv5x_xi302_1505, elementx_x021x_xi300_1479) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi302_1505, elementx_x021x_xi300_1479, tmp_var);
      addx_xi303_1510 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_802_inst
    process(shl92_791, conv95_798) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_791, conv95_798, tmp_var);
      add96_803 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_820_inst
    process(shl98_809, conv101_816) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl98_809, conv101_816, tmp_var);
      add102_821 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_838_inst
    process(shl104_827, conv107_834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl104_827, conv107_834, tmp_var);
      add108_839 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_856_inst
    process(shl110_845, conv113_852) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_845, conv113_852, tmp_var);
      add114_857 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_874_inst
    process(shl116_863, conv119_870) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl116_863, conv119_870, tmp_var);
      add120_875 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_892_inst
    process(shl122_881, conv125_888) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl122_881, conv125_888, tmp_var);
      add126_893 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_910_inst
    process(shl128_899, conv131_906) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl128_899, conv131_906, tmp_var);
      add132_911 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_492_inst
    process(conv9_487) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_487, type_cast_491_wire_constant, tmp_var);
      shl10_493 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_517_inst
    process(conv19_512) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_512, type_cast_516_wire_constant, tmp_var);
      shl20_518 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_542_inst
    process(conv29_537) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_537, type_cast_541_wire_constant, tmp_var);
      shl30_543 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_567_inst
    process(conv39_562) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_562, type_cast_566_wire_constant, tmp_var);
      shl40_568 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_592_inst
    process(conv49_587) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_587, type_cast_591_wire_constant, tmp_var);
      shl50_593 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_617_inst
    process(conv59_612) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_612, type_cast_616_wire_constant, tmp_var);
      shl60_618 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_642_inst
    process(conv69_637) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_637, type_cast_641_wire_constant, tmp_var);
      shl70_643 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_467_inst
    process(conv1_462) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_462, type_cast_466_wire_constant, tmp_var);
      shl_468 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_989_inst
    process(mul82_673) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul82_673, type_cast_988_wire_constant, tmp_var);
      conv2x_xi_990 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1042_inst
    process(addx_xi_1037) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1037, type_cast_1041_wire_constant, tmp_var);
      shl8x_xi_1043 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1069_inst
    process(conv83_679) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv83_679, type_cast_1068_wire_constant, tmp_var);
      Bx_xnot_1070 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1086_inst
    process(shl8x_xix_xlcssa_1060, sh_promx_xi_1082) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xix_xlcssa_1060, sh_promx_xi_1082, tmp_var);
      shl14x_xi_1087 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1136_inst
    process(mul154_1131) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1131, type_cast_1135_wire_constant, tmp_var);
      sext_1137 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1259_inst
    process(conv165_1254) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv165_1254, type_cast_1258_wire_constant, tmp_var);
      shl167_1260 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1277_inst
    process(add171_1272) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_1272, type_cast_1276_wire_constant, tmp_var);
      shl173_1278 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1295_inst
    process(add177_1290) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add177_1290, type_cast_1294_wire_constant, tmp_var);
      shl179_1296 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1313_inst
    process(add183_1308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add183_1308, type_cast_1312_wire_constant, tmp_var);
      shl185_1314 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1331_inst
    process(add189_1326) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add189_1326, type_cast_1330_wire_constant, tmp_var);
      shl191_1332 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1349_inst
    process(add195_1344) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add195_1344, type_cast_1348_wire_constant, tmp_var);
      shl197_1350 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1367_inst
    process(add201_1362) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add201_1362, type_cast_1366_wire_constant, tmp_var);
      shl203_1368 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1414_inst
    process(umax_1409) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1409, type_cast_1413_wire_constant, tmp_var);
      tmp352_1415 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1458_inst
    process(mul154_1131) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1131, type_cast_1457_wire_constant, tmp_var);
      iNsTr_55_1459 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1515_inst
    process(addx_xi303_1510) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi303_1510, type_cast_1514_wire_constant, tmp_var);
      shl8x_xi304_1516 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1542_inst
    process(mul154_1131) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1131, type_cast_1541_wire_constant, tmp_var);
      iNsTr_73_1543 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1559_inst
    process(shl8x_xi304x_xlcssa_1533, sh_promx_xi313_1555) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xi304x_xlcssa_1533, sh_promx_xi313_1555, tmp_var);
      shl14x_xi314_1560 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_790_inst
    process(conv90_785) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv90_785, type_cast_789_wire_constant, tmp_var);
      shl92_791 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_808_inst
    process(add96_803) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add96_803, type_cast_807_wire_constant, tmp_var);
      shl98_809 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_826_inst
    process(add102_821) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add102_821, type_cast_825_wire_constant, tmp_var);
      shl104_827 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_844_inst
    process(add108_839) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_839, type_cast_843_wire_constant, tmp_var);
      shl110_845 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_862_inst
    process(add114_857) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add114_857, type_cast_861_wire_constant, tmp_var);
      shl116_863 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_880_inst
    process(add120_875) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add120_875, type_cast_879_wire_constant, tmp_var);
      shl122_881 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_898_inst
    process(add126_893) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add126_893, type_cast_897_wire_constant, tmp_var);
      shl128_899 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_945_inst
    process(umax365_940) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax365_940, type_cast_944_wire_constant, tmp_var);
      tmp366_946 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1728_inst
    process(conv289_1724, conv230_1716) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv289_1724, conv230_1716, tmp_var);
      sub293_1729 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_684_inst
    process(mul82_673) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_673, type_cast_683_wire_constant, tmp_var);
      cmp325_685 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1151_inst
    process(conv155_1146) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv155_1146, type_cast_1150_wire_constant, tmp_var);
      cmp161321_1152 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1170_inst
    process(tmp350_1165) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp350_1165, type_cast_1169_wire_constant, tmp_var);
      tmp351_1171 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1222_inst
    process(tmp22_1217) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp22_1217, type_cast_1221_wire_constant, tmp_var);
      tmp23_1223 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_718_inst
    process(tmp363_713) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp363_713, type_cast_717_wire_constant, tmp_var);
      tmp364_719 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_753_inst
    process(tmp30_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp30_748, type_cast_752_wire_constant, tmp_var);
      tmp31_754 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1051_inst
    process(convx_xi_1047, shlx_xi_996) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_1047, shlx_xi_996, tmp_var);
      cmpx_xi_1052 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1524_inst
    process(convx_xi305_1520, shlx_xi297_1469) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi305_1520, shlx_xi297_1469, tmp_var);
      cmpx_xi306_1525 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1081_inst
    process(add1216x_xi_1076) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi_1076, type_cast_1080_wire_constant, tmp_var);
      sh_promx_xi_1082 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1554_inst
    process(add1216x_xi312_1549) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi312_1549, type_cast_1553_wire_constant, tmp_var);
      sh_promx_xi313_1555 <= tmp_var; --
    end process;
    -- shared split operator group (116) : array_obj_ref_1092_index_offset 
    ApIntAdd_group_116: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1091_scaled;
      array_obj_ref_1092_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1092_index_offset_req_0;
      array_obj_ref_1092_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1092_index_offset_req_1;
      array_obj_ref_1092_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_116_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_116_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_116",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 116
    -- shared split operator group (117) : array_obj_ref_1245_index_offset 
    ApIntAdd_group_117: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar355_1244_scaled;
      array_obj_ref_1245_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1245_index_offset_req_0;
      array_obj_ref_1245_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1245_index_offset_req_1;
      array_obj_ref_1245_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_117_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_117_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- shared split operator group (118) : array_obj_ref_1565_index_offset 
    ApIntAdd_group_118: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_1564_scaled;
      array_obj_ref_1565_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1565_index_offset_req_0;
      array_obj_ref_1565_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1565_index_offset_req_1;
      array_obj_ref_1565_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_118_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_118_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- shared split operator group (119) : array_obj_ref_776_index_offset 
    ApIntAdd_group_119: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar369_775_scaled;
      array_obj_ref_776_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_776_index_offset_req_0;
      array_obj_ref_776_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_776_index_offset_req_1;
      array_obj_ref_776_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_119_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_119_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_119",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 119
    -- unary operator type_cast_1209_inst
    process(tmp20_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp20_1206, tmp_var);
      type_cast_1209_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1714_inst
    process(call229_1576) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call229_1576, tmp_var);
      type_cast_1714_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1722_inst
    process(call288_1719) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call288_1719, tmp_var);
      type_cast_1722_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_677_inst
    process(mul82_673) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul82_673, tmp_var);
      type_cast_677_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_705_inst
    process(tmp361_702) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp361_702, tmp_var);
      type_cast_705_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_740_inst
    process(tmp28_737) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp28_737, tmp_var);
      type_cast_740_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_913_store_0 ptr_deref_1096_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_913_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1096_store_0_req_0;
      ptr_deref_913_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1096_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_913_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1096_store_0_req_1;
      ptr_deref_913_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1096_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_913_word_address_0 & ptr_deref_1096_word_address_0;
      data_in <= ptr_deref_913_data_0 & ptr_deref_1096_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1382_store_0 ptr_deref_1569_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1382_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1569_store_0_req_0;
      ptr_deref_1382_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1569_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1382_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1569_store_0_req_1;
      ptr_deref_1382_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1569_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1382_word_address_0 & ptr_deref_1569_word_address_0;
      data_in <= ptr_deref_1382_data_0 & ptr_deref_1569_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_570_inst RPIPE_maxpool_input_pipe_470_inst RPIPE_maxpool_input_pipe_545_inst RPIPE_maxpool_input_pipe_482_inst RPIPE_maxpool_input_pipe_620_inst RPIPE_maxpool_input_pipe_495_inst RPIPE_maxpool_input_pipe_557_inst RPIPE_maxpool_input_pipe_645_inst RPIPE_maxpool_input_pipe_507_inst RPIPE_maxpool_input_pipe_595_inst RPIPE_maxpool_input_pipe_582_inst RPIPE_maxpool_input_pipe_632_inst RPIPE_maxpool_input_pipe_520_inst RPIPE_maxpool_input_pipe_532_inst RPIPE_maxpool_input_pipe_607_inst RPIPE_maxpool_input_pipe_847_inst RPIPE_maxpool_input_pipe_1027_inst RPIPE_maxpool_input_pipe_793_inst RPIPE_maxpool_input_pipe_901_inst RPIPE_maxpool_input_pipe_811_inst RPIPE_maxpool_input_pipe_883_inst RPIPE_maxpool_input_pipe_865_inst RPIPE_maxpool_input_pipe_780_inst RPIPE_maxpool_input_pipe_829_inst RPIPE_maxpool_input_pipe_457_inst RPIPE_maxpool_input_pipe_1249_inst RPIPE_maxpool_input_pipe_1262_inst RPIPE_maxpool_input_pipe_1280_inst RPIPE_maxpool_input_pipe_1298_inst RPIPE_maxpool_input_pipe_1316_inst RPIPE_maxpool_input_pipe_1334_inst RPIPE_maxpool_input_pipe_1352_inst RPIPE_maxpool_input_pipe_1370_inst RPIPE_maxpool_input_pipe_1500_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_570_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_470_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_545_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_482_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_620_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_495_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_557_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_645_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_507_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_595_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_582_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_632_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_520_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_532_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_607_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_847_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_1027_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_793_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_901_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_811_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_883_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_865_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_780_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_829_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_457_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_1249_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_1262_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_1280_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_1298_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_1316_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_1334_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_1352_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1370_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1500_inst_req_0;
      RPIPE_maxpool_input_pipe_570_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_470_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_545_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_482_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_620_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_495_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_557_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_645_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_507_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_595_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_582_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_632_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_520_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_532_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_607_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_847_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_1027_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_793_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_901_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_811_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_883_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_865_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_780_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_829_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_457_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_1249_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_1262_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_1280_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_1298_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_1316_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_1334_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_1352_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1370_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1500_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_570_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_470_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_545_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_482_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_620_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_495_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_557_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_645_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_507_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_595_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_582_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_632_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_520_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_532_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_607_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_847_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_1027_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_793_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_901_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_811_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_883_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_865_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_780_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_829_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_457_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_1249_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_1262_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_1280_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_1298_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_1316_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_1334_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_1352_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1370_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1500_inst_req_1;
      RPIPE_maxpool_input_pipe_570_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_470_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_545_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_482_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_620_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_495_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_557_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_645_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_507_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_595_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_582_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_632_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_520_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_532_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_607_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_847_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_1027_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_793_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_901_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_811_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_883_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_865_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_780_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_829_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_457_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_1249_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_1262_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_1280_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_1298_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_1316_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_1334_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_1352_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1370_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1500_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call41_571 <= data_out(271 downto 264);
      call2_471 <= data_out(263 downto 256);
      call31_546 <= data_out(255 downto 248);
      call6_483 <= data_out(247 downto 240);
      call61_621 <= data_out(239 downto 232);
      call11_496 <= data_out(231 downto 224);
      call36_558 <= data_out(223 downto 216);
      call71_646 <= data_out(215 downto 208);
      call16_508 <= data_out(207 downto 200);
      call51_596 <= data_out(199 downto 192);
      call46_583 <= data_out(191 downto 184);
      call66_633 <= data_out(183 downto 176);
      call21_521 <= data_out(175 downto 168);
      call26_533 <= data_out(167 downto 160);
      call56_608 <= data_out(159 downto 152);
      call111_848 <= data_out(151 downto 144);
      callx_xi_1028 <= data_out(143 downto 136);
      call93_794 <= data_out(135 downto 128);
      call129_902 <= data_out(127 downto 120);
      call99_812 <= data_out(119 downto 112);
      call123_884 <= data_out(111 downto 104);
      call117_866 <= data_out(103 downto 96);
      call89_781 <= data_out(95 downto 88);
      call105_830 <= data_out(87 downto 80);
      call_458 <= data_out(79 downto 72);
      call164_1250 <= data_out(71 downto 64);
      call168_1263 <= data_out(63 downto 56);
      call174_1281 <= data_out(55 downto 48);
      call180_1299 <= data_out(47 downto 40);
      call186_1317 <= data_out(39 downto 32);
      call192_1335 <= data_out(31 downto 24);
      call198_1353 <= data_out(23 downto 16);
      call204_1371 <= data_out(15 downto 8);
      callx_xi301_1501 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_1730_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1730_inst_req_0;
      WPIPE_elapsed_time_pipe_1730_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1730_inst_req_1;
      WPIPE_elapsed_time_pipe_1730_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub293_1729;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_maxpool_output_pipe_1583_inst WPIPE_maxpool_output_pipe_1587_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1583_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1587_inst_req_0;
      WPIPE_maxpool_output_pipe_1583_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1587_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1583_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1587_inst_req_1;
      WPIPE_maxpool_output_pipe_1583_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1587_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= type_cast_1585_wire_constant & type_cast_1589_wire_constant;
      maxpool_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_num_out_pipe_1666_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_1666_inst_req_0;
      WPIPE_num_out_pipe_1666_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_num_out_pipe_1666_inst_req_1;
      WPIPE_num_out_pipe_1666_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= mul249_1595;
      num_out_pipe_write_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_1576_call call_stmt_1719_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1576_call_req_0;
      reqL_unguarded(0) <= call_stmt_1719_call_req_0;
      call_stmt_1576_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1719_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1576_call_req_1;
      reqR_unguarded(0) <= call_stmt_1719_call_req_1;
      call_stmt_1576_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1719_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call229_1576 <= data_out(127 downto 64);
      call288_1719 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1686_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(135 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1686_call_req_0;
      call_stmt_1686_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1686_call_req_1;
      call_stmt_1686_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv255_1672 & conv261_1676 & and264_1682;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 136,
        owidth => 136,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(135 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1693_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1693_call_req_0;
      call_stmt_1693_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1693_call_req_1;
      call_stmt_1693_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul236_1582 & add33_555 & sub_1601 & sub273_1607 & add23_530 & add13_505;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 96,
        owidth => 96,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(95 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_3851_start: Boolean;
  signal convolve_CP_3851_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_1766_ack_0 : boolean;
  signal nmycount_1840_1768_buf_ack_1 : boolean;
  signal nacc_1832_1772_buf_req_1 : boolean;
  signal nmycount_1840_1768_buf_req_1 : boolean;
  signal phi_stmt_1774_req_1 : boolean;
  signal do_while_stmt_1764_branch_req_0 : boolean;
  signal nacc_1832_1772_buf_req_0 : boolean;
  signal phi_stmt_1774_ack_0 : boolean;
  signal slice_1753_inst_req_1 : boolean;
  signal phi_stmt_1774_req_0 : boolean;
  signal slice_1753_inst_ack_1 : boolean;
  signal nacc_1832_1772_buf_ack_1 : boolean;
  signal phi_stmt_1770_req_0 : boolean;
  signal phi_stmt_1770_req_1 : boolean;
  signal nacc_1832_1772_buf_ack_0 : boolean;
  signal phi_stmt_1766_req_0 : boolean;
  signal nmycount_1840_1768_buf_req_0 : boolean;
  signal nmycount_1840_1768_buf_ack_0 : boolean;
  signal phi_stmt_1766_req_1 : boolean;
  signal phi_stmt_1770_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1742_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1742_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1742_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1742_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_1745_inst_req_0 : boolean;
  signal RPIPE_size_pipe_1745_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_1745_inst_req_1 : boolean;
  signal RPIPE_size_pipe_1745_inst_ack_1 : boolean;
  signal slice_1749_inst_req_0 : boolean;
  signal slice_1749_inst_ack_0 : boolean;
  signal slice_1749_inst_req_1 : boolean;
  signal slice_1749_inst_ack_1 : boolean;
  signal slice_1753_inst_req_0 : boolean;
  signal slice_1753_inst_ack_0 : boolean;
  signal n_out_count_1881_1778_buf_req_0 : boolean;
  signal n_out_count_1881_1778_buf_ack_0 : boolean;
  signal n_out_count_1881_1778_buf_req_1 : boolean;
  signal n_out_count_1881_1778_buf_ack_1 : boolean;
  signal RPIPE_input_pipe1_1781_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_1781_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_1781_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_1781_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_1789_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe1_1789_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_1789_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_1789_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe2_1793_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe2_1793_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe2_1793_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe2_1793_inst_ack_1 : boolean;
  signal SUB_u31_u31_1813_inst_req_0 : boolean;
  signal SUB_u31_u31_1813_inst_ack_0 : boolean;
  signal SUB_u31_u31_1813_inst_req_1 : boolean;
  signal SUB_u31_u31_1813_inst_ack_1 : boolean;
  signal NOT_u1_u1_1848_inst_req_0 : boolean;
  signal NOT_u1_u1_1848_inst_ack_0 : boolean;
  signal NOT_u1_u1_1848_inst_req_1 : boolean;
  signal NOT_u1_u1_1848_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_1863_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_1863_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_1863_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_1863_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe2_1867_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_1867_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_1867_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe2_1867_inst_ack_1 : boolean;
  signal WPIPE_input_done_pipe_1888_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_1888_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_1888_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_1888_inst_ack_1 : boolean;
  signal slice_1893_inst_req_0 : boolean;
  signal slice_1893_inst_ack_0 : boolean;
  signal slice_1893_inst_req_1 : boolean;
  signal slice_1893_inst_ack_1 : boolean;
  signal slice_1897_inst_req_0 : boolean;
  signal slice_1897_inst_ack_0 : boolean;
  signal slice_1897_inst_req_1 : boolean;
  signal slice_1897_inst_ack_1 : boolean;
  signal W_next_sum_1872_delayed_1_0_1899_inst_req_0 : boolean;
  signal W_next_sum_1872_delayed_1_0_1899_inst_ack_0 : boolean;
  signal W_next_sum_1872_delayed_1_0_1899_inst_req_1 : boolean;
  signal W_next_sum_1872_delayed_1_0_1899_inst_ack_1 : boolean;
  signal type_cast_1905_inst_req_0 : boolean;
  signal type_cast_1905_inst_ack_0 : boolean;
  signal type_cast_1905_inst_req_1 : boolean;
  signal type_cast_1905_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1903_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1903_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1903_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1903_inst_ack_1 : boolean;
  signal W_next_sum_1877_delayed_1_0_1907_inst_req_0 : boolean;
  signal W_next_sum_1877_delayed_1_0_1907_inst_ack_0 : boolean;
  signal W_next_sum_1877_delayed_1_0_1907_inst_req_1 : boolean;
  signal W_next_sum_1877_delayed_1_0_1907_inst_ack_1 : boolean;
  signal type_cast_1913_inst_req_0 : boolean;
  signal type_cast_1913_inst_ack_0 : boolean;
  signal type_cast_1913_inst_req_1 : boolean;
  signal type_cast_1913_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1911_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1911_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1911_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1911_inst_ack_1 : boolean;
  signal do_while_stmt_1764_branch_ack_0 : boolean;
  signal do_while_stmt_1764_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_3851_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_3851_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_3851_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_3851_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_3851: Block -- control-path 
    signal convolve_CP_3851_elements: BooleanArray(144 downto 0);
    -- 
  begin -- 
    convolve_CP_3851_elements(0) <= convolve_CP_3851_start;
    convolve_CP_3851_symbol <= convolve_CP_3851_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	144 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1739/$entry
      -- CP-element group 0: 	 branch_block_stmt_1739/branch_block_stmt_1739__entry__
      -- CP-element group 0: 	 branch_block_stmt_1739/merge_stmt_1740__entry__
      -- CP-element group 0: 	 branch_block_stmt_1739/merge_stmt_1740_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1739/merge_stmt_1740__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1739/merge_stmt_1740__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1739/$exit
      -- CP-element group 1: 	 branch_block_stmt_1739/branch_block_stmt_1739__exit__
      -- 
    convolve_CP_3851_elements(1) <= false; 
    -- CP-element group 2:  transition  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	143 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	144 
    -- CP-element group 2:  members (4) 
      -- CP-element group 2: 	 branch_block_stmt_1739/do_while_stmt_1764__exit__
      -- CP-element group 2: 	 branch_block_stmt_1739/loopback
      -- CP-element group 2: 	 branch_block_stmt_1739/loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1739/loopback_PhiReq/$exit
      -- 
    convolve_CP_3851_elements(2) <= convolve_CP_3851_elements(143);
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	144 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_Update/cr
      -- 
    ra_3877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1742_inst_ack_0, ack => convolve_CP_3851_elements(3)); -- 
    cr_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(3), ack => RPIPE_num_out_pipe_1742_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	11 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_Update/ca
      -- 
    ca_3882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1742_inst_ack_1, ack => convolve_CP_3851_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	144 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_Update/cr
      -- 
    ra_3891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1745_inst_ack_0, ack => convolve_CP_3851_elements(5)); -- 
    cr_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(5), ack => RPIPE_size_pipe_1745_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_Sample/rr
      -- 
    ca_3896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1745_inst_ack_1, ack => convolve_CP_3851_elements(6)); -- 
    rr_3904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(6), ack => slice_1749_inst_req_0); -- 
    rr_3918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(6), ack => slice_1753_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_Sample/ra
      -- 
    ra_3905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1749_inst_ack_0, ack => convolve_CP_3851_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	144 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_Update/ca
      -- 
    ca_3910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1749_inst_ack_1, ack => convolve_CP_3851_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_Sample/ra
      -- 
    ra_3919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1753_inst_ack_0, ack => convolve_CP_3851_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	144 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_update_completed_
      -- 
    ca_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1753_inst_ack_1, ack => convolve_CP_3851_elements(10)); -- 
    -- CP-element group 11:  join  transition  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: 	4 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763__exit__
      -- CP-element group 11: 	 branch_block_stmt_1739/do_while_stmt_1764__entry__
      -- CP-element group 11: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/$exit
      -- 
    convolve_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(10) & convolve_CP_3851_elements(4) & convolve_CP_3851_elements(8);
      gj_convolve_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	18 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764__entry__
      -- CP-element group 12: 	 branch_block_stmt_1739/do_while_stmt_1764/$entry
      -- 
    convolve_CP_3851_elements(12) <= convolve_CP_3851_elements(11);
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	143 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764__exit__
      -- 
    -- Element group convolve_CP_3851_elements(13) is bound as output of CP function.
    -- CP-element group 14:  merge  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1739/do_while_stmt_1764/loop_back
      -- 
    -- Element group convolve_CP_3851_elements(14) is bound as output of CP function.
    -- CP-element group 15:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	141 
    -- CP-element group 15: 	142 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1739/do_while_stmt_1764/condition_done
      -- CP-element group 15: 	 branch_block_stmt_1739/do_while_stmt_1764/loop_exit/$entry
      -- CP-element group 15: 	 branch_block_stmt_1739/do_while_stmt_1764/loop_taken/$entry
      -- 
    convolve_CP_3851_elements(15) <= convolve_CP_3851_elements(20);
    -- CP-element group 16:  branch  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	140 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1739/do_while_stmt_1764/loop_body_done
      -- 
    convolve_CP_3851_elements(16) <= convolve_CP_3851_elements(140);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	67 
    -- CP-element group 17: 	50 
    -- CP-element group 17: 	31 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_3851_elements(17) <= convolve_CP_3851_elements(14);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	12 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	69 
    -- CP-element group 18: 	52 
    -- CP-element group 18: 	33 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_3851_elements(18) <= convolve_CP_3851_elements(12);
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	139 
    -- CP-element group 19: 	25 
    -- CP-element group 19: 	26 
    -- CP-element group 19: 	80 
    -- CP-element group 19: 	84 
    -- CP-element group 19: 	88 
    -- CP-element group 19: 	92 
    -- CP-element group 19: 	63 
    -- CP-element group 19: 	64 
    -- CP-element group 19: 	96 
    -- CP-element group 19: 	44 
    -- CP-element group 19: 	45 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/loop_body_start
      -- CP-element group 19: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/$entry
      -- 
    -- Element group convolve_CP_3851_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	139 
    -- CP-element group 20: 	66 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	95 
    -- CP-element group 20: 	30 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/condition_evaluated
      -- 
    condition_evaluated_3939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(20), ack => do_while_stmt_1764_branch_req_0); -- 
    convolve_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(139) & convolve_CP_3851_elements(66) & convolve_CP_3851_elements(24) & convolve_CP_3851_elements(95) & convolve_CP_3851_elements(30);
      gj_convolve_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	25 
    -- CP-element group 21: 	63 
    -- CP-element group 21: 	44 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	27 
    -- CP-element group 21: 	46 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/aggregated_phi_sample_req
      -- CP-element group 21: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_sample_start__ps
      -- 
    convolve_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(25) & convolve_CP_3851_elements(63) & convolve_CP_3851_elements(44) & convolve_CP_3851_elements(24);
      gj_convolve_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	65 
    -- CP-element group 22: 	47 
    -- CP-element group 22: 	28 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	81 
    -- CP-element group 22: 	85 
    -- CP-element group 22: 	89 
    -- CP-element group 22: 	93 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	63 
    -- CP-element group 22: 	44 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/aggregated_phi_sample_ack
      -- CP-element group 22: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_sample_completed_
      -- 
    convolve_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(65) & convolve_CP_3851_elements(47) & convolve_CP_3851_elements(28);
      gj_convolve_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	26 
    -- CP-element group 23: 	64 
    -- CP-element group 23: 	45 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	48 
    -- CP-element group 23: 	29 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_update_start__ps
      -- CP-element group 23: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/aggregated_phi_update_req
      -- 
    convolve_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(26) & convolve_CP_3851_elements(64) & convolve_CP_3851_elements(45);
      gj_convolve_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	66 
    -- CP-element group 24: 	49 
    -- CP-element group 24: 	30 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	21 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(66) & convolve_CP_3851_elements(49) & convolve_CP_3851_elements(30);
      gj_convolve_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	19 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	95 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	21 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_sample_start_
      -- 
    convolve_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(95) & convolve_CP_3851_elements(22);
      gj_convolve_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	19 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	119 
    -- CP-element group 26: 	130 
    -- CP-element group 26: 	30 
    -- CP-element group 26: 	107 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	23 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_update_start_
      -- 
    convolve_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(119) & convolve_CP_3851_elements(130) & convolve_CP_3851_elements(30) & convolve_CP_3851_elements(107);
      gj_convolve_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	21 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_sample_start__ps
      -- 
    convolve_CP_3851_elements(27) <= convolve_CP_3851_elements(21);
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	22 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_sample_completed__ps
      -- 
    -- Element group convolve_CP_3851_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_update_start__ps
      -- 
    convolve_CP_3851_elements(29) <= convolve_CP_3851_elements(23);
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: 	117 
    -- CP-element group 30: 	106 
    -- CP-element group 30: 	128 
    -- CP-element group 30: 	20 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	26 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_update_completed__ps
      -- 
    -- Element group convolve_CP_3851_elements(30) is bound as output of CP function.
    -- CP-element group 31:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	17 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_loopback_trigger
      -- 
    convolve_CP_3851_elements(31) <= convolve_CP_3851_elements(17);
    -- CP-element group 32:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_loopback_sample_req
      -- CP-element group 32: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_loopback_sample_req_ps
      -- 
    phi_stmt_1766_loopback_sample_req_3954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1766_loopback_sample_req_3954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(32), ack => phi_stmt_1766_req_0); -- 
    -- Element group convolve_CP_3851_elements(32) is bound as output of CP function.
    -- CP-element group 33:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	18 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_entry_trigger
      -- 
    convolve_CP_3851_elements(33) <= convolve_CP_3851_elements(18);
    -- CP-element group 34:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_entry_sample_req_ps
      -- CP-element group 34: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_entry_sample_req
      -- 
    phi_stmt_1766_entry_sample_req_3957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1766_entry_sample_req_3957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(34), ack => phi_stmt_1766_req_1); -- 
    -- Element group convolve_CP_3851_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_phi_mux_ack
      -- CP-element group 35: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1766_phi_mux_ack_ps
      -- 
    phi_stmt_1766_phi_mux_ack_3960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1766_ack_0, ack => convolve_CP_3851_elements(35)); -- 
    -- CP-element group 36:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_sample_start__ps
      -- CP-element group 36: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_Sample/req
      -- 
    req_3973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(36), ack => nmycount_1840_1768_buf_req_0); -- 
    -- Element group convolve_CP_3851_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_Update/req
      -- CP-element group 37: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_update_start__ps
      -- CP-element group 37: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_update_start_
      -- 
    req_3978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(37), ack => nmycount_1840_1768_buf_req_1); -- 
    -- Element group convolve_CP_3851_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_sample_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_Sample/ack
      -- 
    ack_3974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1840_1768_buf_ack_0, ack => convolve_CP_3851_elements(38)); -- 
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_update_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nmycount_1768_update_completed_
      -- 
    ack_3979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1840_1768_buf_ack_1, ack => convolve_CP_3851_elements(39)); -- 
    -- CP-element group 40:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_mcount_var_1769_sample_start__ps
      -- CP-element group 40: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_mcount_var_1769_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_mcount_var_1769_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_mcount_var_1769_sample_completed__ps
      -- 
    -- Element group convolve_CP_3851_elements(40) is bound as output of CP function.
    -- CP-element group 41:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_mcount_var_1769_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_mcount_var_1769_update_start__ps
      -- 
    -- Element group convolve_CP_3851_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_mcount_var_1769_update_completed__ps
      -- 
    convolve_CP_3851_elements(42) <= convolve_CP_3851_elements(43);
    -- CP-element group 43:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	42 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_mcount_var_1769_update_completed_
      -- 
    -- Element group convolve_CP_3851_elements(43) is a control-delay.
    cp_element_43_delay: control_delay_element  generic map(name => " 43_delay", delay_value => 1)  port map(req => convolve_CP_3851_elements(41), ack => convolve_CP_3851_elements(43), clk => clk, reset =>reset);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	19 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	83 
    -- CP-element group 44: 	87 
    -- CP-element group 44: 	91 
    -- CP-element group 44: 	95 
    -- CP-element group 44: 	22 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_sample_start_
      -- 
    convolve_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(83) & convolve_CP_3851_elements(87) & convolve_CP_3851_elements(91) & convolve_CP_3851_elements(95) & convolve_CP_3851_elements(22);
      gj_convolve_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	19 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	49 
    -- CP-element group 45: 	115 
    -- CP-element group 45: 	111 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	23 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_update_start_
      -- 
    convolve_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(49) & convolve_CP_3851_elements(115) & convolve_CP_3851_elements(111);
      gj_convolve_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	21 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_sample_start__ps
      -- 
    convolve_CP_3851_elements(46) <= convolve_CP_3851_elements(21);
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	22 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_sample_completed__ps
      -- 
    -- Element group convolve_CP_3851_elements(47) is bound as output of CP function.
    -- CP-element group 48:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	23 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_update_start__ps
      -- 
    convolve_CP_3851_elements(48) <= convolve_CP_3851_elements(23);
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	24 
    -- CP-element group 49: 	113 
    -- CP-element group 49: 	109 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	45 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_update_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_update_completed_
      -- 
    -- Element group convolve_CP_3851_elements(49) is bound as output of CP function.
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	17 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_loopback_trigger
      -- 
    convolve_CP_3851_elements(50) <= convolve_CP_3851_elements(17);
    -- CP-element group 51:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_loopback_sample_req
      -- CP-element group 51: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_loopback_sample_req_ps
      -- 
    phi_stmt_1770_loopback_sample_req_3998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1770_loopback_sample_req_3998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(51), ack => phi_stmt_1770_req_0); -- 
    -- Element group convolve_CP_3851_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	18 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_entry_trigger
      -- 
    convolve_CP_3851_elements(52) <= convolve_CP_3851_elements(18);
    -- CP-element group 53:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_entry_sample_req_ps
      -- CP-element group 53: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_entry_sample_req
      -- 
    phi_stmt_1770_entry_sample_req_4001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1770_entry_sample_req_4001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(53), ack => phi_stmt_1770_req_1); -- 
    -- Element group convolve_CP_3851_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_phi_mux_ack_ps
      -- CP-element group 54: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1770_phi_mux_ack
      -- 
    phi_stmt_1770_phi_mux_ack_4004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1770_ack_0, ack => convolve_CP_3851_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_sample_start__ps
      -- CP-element group 55: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_Sample/req
      -- CP-element group 55: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_sample_start_
      -- 
    req_4017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(55), ack => nacc_1832_1772_buf_req_0); -- 
    -- Element group convolve_CP_3851_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_Update/req
      -- CP-element group 56: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_update_start_
      -- CP-element group 56: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_update_start__ps
      -- CP-element group 56: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_Update/$entry
      -- 
    req_4022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(56), ack => nacc_1832_1772_buf_req_1); -- 
    -- Element group convolve_CP_3851_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_sample_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_sample_completed_
      -- 
    ack_4018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1832_1772_buf_ack_0, ack => convolve_CP_3851_elements(57)); -- 
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_update_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_nacc_1772_Update/$exit
      -- 
    ack_4023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1832_1772_buf_ack_1, ack => convolve_CP_3851_elements(58)); -- 
    -- CP-element group 59:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_acc_var_1773_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_acc_var_1773_sample_start__ps
      -- CP-element group 59: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_acc_var_1773_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_acc_var_1773_sample_completed__ps
      -- 
    -- Element group convolve_CP_3851_elements(59) is bound as output of CP function.
    -- CP-element group 60:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_acc_var_1773_update_start__ps
      -- CP-element group 60: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_acc_var_1773_update_start_
      -- 
    -- Element group convolve_CP_3851_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_acc_var_1773_update_completed__ps
      -- 
    convolve_CP_3851_elements(61) <= convolve_CP_3851_elements(62);
    -- CP-element group 62:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	61 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_acc_var_1773_update_completed_
      -- 
    -- Element group convolve_CP_3851_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => convolve_CP_3851_elements(60), ack => convolve_CP_3851_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  join  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	19 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	95 
    -- CP-element group 63: 	22 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	21 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_sample_start_
      -- 
    convolve_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(95) & convolve_CP_3851_elements(22);
      gj_convolve_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	19 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: 	101 
    -- CP-element group 64: 	104 
    -- CP-element group 64: 	107 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	23 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_update_start_
      -- 
    convolve_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(66) & convolve_CP_3851_elements(101) & convolve_CP_3851_elements(104) & convolve_CP_3851_elements(107);
      gj_convolve_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	22 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_sample_completed__ps
      -- 
    -- Element group convolve_CP_3851_elements(65) is bound as output of CP function.
    -- CP-element group 66:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	24 
    -- CP-element group 66: 	103 
    -- CP-element group 66: 	106 
    -- CP-element group 66: 	100 
    -- CP-element group 66: 	20 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_update_completed__ps
      -- 
    -- Element group convolve_CP_3851_elements(66) is bound as output of CP function.
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	17 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_loopback_trigger
      -- 
    convolve_CP_3851_elements(67) <= convolve_CP_3851_elements(17);
    -- CP-element group 68:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_loopback_sample_req
      -- CP-element group 68: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_loopback_sample_req_ps
      -- 
    phi_stmt_1774_loopback_sample_req_4042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1774_loopback_sample_req_4042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(68), ack => phi_stmt_1774_req_1); -- 
    -- Element group convolve_CP_3851_elements(68) is bound as output of CP function.
    -- CP-element group 69:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	18 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_entry_trigger
      -- 
    convolve_CP_3851_elements(69) <= convolve_CP_3851_elements(18);
    -- CP-element group 70:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_entry_sample_req
      -- CP-element group 70: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_entry_sample_req_ps
      -- 
    phi_stmt_1774_entry_sample_req_4045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1774_entry_sample_req_4045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(70), ack => phi_stmt_1774_req_0); -- 
    -- Element group convolve_CP_3851_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_phi_mux_ack
      -- CP-element group 71: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/phi_stmt_1774_phi_mux_ack_ps
      -- 
    phi_stmt_1774_phi_mux_ack_4048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1774_ack_0, ack => convolve_CP_3851_elements(71)); -- 
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1777_sample_completed__ps
      -- CP-element group 72: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1777_sample_start__ps
      -- CP-element group 72: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1777_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1777_sample_completed_
      -- 
    -- Element group convolve_CP_3851_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1777_update_start_
      -- CP-element group 73: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1777_update_start__ps
      -- 
    -- Element group convolve_CP_3851_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1777_update_completed__ps
      -- 
    convolve_CP_3851_elements(74) <= convolve_CP_3851_elements(75);
    -- CP-element group 75:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	74 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1777_update_completed_
      -- 
    -- Element group convolve_CP_3851_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convolve_CP_3851_elements(73), ack => convolve_CP_3851_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_sample_start__ps
      -- CP-element group 76: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_Sample/req
      -- 
    req_4069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(76), ack => n_out_count_1881_1778_buf_req_0); -- 
    -- Element group convolve_CP_3851_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_update_start__ps
      -- CP-element group 77: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_Update/req
      -- 
    req_4074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(77), ack => n_out_count_1881_1778_buf_req_1); -- 
    -- Element group convolve_CP_3851_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (4) 
      -- CP-element group 78: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_sample_completed__ps
      -- CP-element group 78: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_Sample/ack
      -- 
    ack_4070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1881_1778_buf_ack_0, ack => convolve_CP_3851_elements(78)); -- 
    -- CP-element group 79:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_update_completed__ps
      -- CP-element group 79: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/R_n_out_count_1778_Update/ack
      -- 
    ack_4075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1881_1778_buf_ack_1, ack => convolve_CP_3851_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	19 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	83 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_Sample/rr
      -- 
    rr_4084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(80), ack => RPIPE_input_pipe1_1781_inst_req_0); -- 
    convolve_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(83);
      gj_convolve_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: 	22 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	115 
    -- CP-element group 81: 	111 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_Update/cr
      -- 
    cr_4089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(81), ack => RPIPE_input_pipe1_1781_inst_req_1); -- 
    convolve_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(82) & convolve_CP_3851_elements(22) & convolve_CP_3851_elements(115) & convolve_CP_3851_elements(111);
      gj_convolve_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	81 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_Sample/ra
      -- 
    ra_4085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1781_inst_ack_0, ack => convolve_CP_3851_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	113 
    -- CP-element group 83: 	109 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	44 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_input_pipe1_1781_Update/ca
      -- 
    ca_4090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1781_inst_ack_1, ack => convolve_CP_3851_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	19 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	87 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_Sample/rr
      -- 
    rr_4098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(84), ack => RPIPE_kernel_pipe1_1789_inst_req_0); -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(87);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: 	22 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	115 
    -- CP-element group 85: 	101 
    -- CP-element group 85: 	104 
    -- CP-element group 85: 	111 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_Update/cr
      -- 
    cr_4103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(85), ack => RPIPE_kernel_pipe1_1789_inst_req_1); -- 
    convolve_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 15,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(86) & convolve_CP_3851_elements(22) & convolve_CP_3851_elements(115) & convolve_CP_3851_elements(101) & convolve_CP_3851_elements(104) & convolve_CP_3851_elements(111);
      gj_convolve_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	85 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_Sample/ra
      -- 
    ra_4099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1789_inst_ack_0, ack => convolve_CP_3851_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	113 
    -- CP-element group 87: 	103 
    -- CP-element group 87: 	100 
    -- CP-element group 87: 	109 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	84 
    -- CP-element group 87: 	44 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe1_1789_Update/ca
      -- 
    ca_4104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1789_inst_ack_1, ack => convolve_CP_3851_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	19 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	91 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_Sample/rr
      -- 
    rr_4112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(88), ack => RPIPE_kernel_pipe2_1793_inst_req_0); -- 
    convolve_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(91);
      gj_convolve_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	22 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	115 
    -- CP-element group 89: 	101 
    -- CP-element group 89: 	104 
    -- CP-element group 89: 	111 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_Update/cr
      -- 
    cr_4117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(89), ack => RPIPE_kernel_pipe2_1793_inst_req_1); -- 
    convolve_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 15,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(90) & convolve_CP_3851_elements(22) & convolve_CP_3851_elements(115) & convolve_CP_3851_elements(101) & convolve_CP_3851_elements(104) & convolve_CP_3851_elements(111);
      gj_convolve_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_Sample/ra
      -- 
    ra_4113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_1793_inst_ack_0, ack => convolve_CP_3851_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	113 
    -- CP-element group 91: 	103 
    -- CP-element group 91: 	100 
    -- CP-element group 91: 	109 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	88 
    -- CP-element group 91: 	44 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/RPIPE_kernel_pipe2_1793_Update/ca
      -- 
    ca_4118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_1793_inst_ack_1, ack => convolve_CP_3851_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	19 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_Sample/rr
      -- 
    rr_4126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(92), ack => SUB_u31_u31_1813_inst_req_0); -- 
    convolve_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(94);
      gj_convolve_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	22 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	119 
    -- CP-element group 93: 	130 
    -- CP-element group 93: 	95 
    -- CP-element group 93: 	107 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_update_start_
      -- CP-element group 93: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_Update/cr
      -- 
    cr_4131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(93), ack => SUB_u31_u31_1813_inst_req_1); -- 
    convolve_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(22) & convolve_CP_3851_elements(119) & convolve_CP_3851_elements(130) & convolve_CP_3851_elements(95) & convolve_CP_3851_elements(107);
      gj_convolve_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_Sample/ra
      -- 
    ra_4127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u31_u31_1813_inst_ack_0, ack => convolve_CP_3851_elements(94)); -- 
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	117 
    -- CP-element group 95: 	106 
    -- CP-element group 95: 	128 
    -- CP-element group 95: 	20 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	25 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	63 
    -- CP-element group 95: 	44 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/SUB_u31_u31_1813_Update/ca
      -- 
    ca_4132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u31_u31_1813_inst_ack_1, ack => convolve_CP_3851_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	19 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_Sample/rr
      -- 
    rr_4140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(96), ack => NOT_u1_u1_1848_inst_req_0); -- 
    convolve_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(19) & convolve_CP_3851_elements(98);
      gj_convolve_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	101 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_update_start_
      -- CP-element group 97: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_Update/cr
      -- 
    cr_4145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(97), ack => NOT_u1_u1_1848_inst_req_1); -- 
    convolve_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(101) & convolve_CP_3851_elements(99);
      gj_convolve_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_Sample/ra
      -- 
    ra_4141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1848_inst_ack_0, ack => convolve_CP_3851_elements(98)); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/NOT_u1_u1_1848_Update/ca
      -- 
    ca_4146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1848_inst_ack_1, ack => convolve_CP_3851_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	66 
    -- CP-element group 100: 	87 
    -- CP-element group 100: 	91 
    -- CP-element group 100: 	99 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_Sample/req
      -- 
    req_4154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(100), ack => WPIPE_kernel_pipe1_1863_inst_req_0); -- 
    convolve_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(66) & convolve_CP_3851_elements(87) & convolve_CP_3851_elements(91) & convolve_CP_3851_elements(99) & convolve_CP_3851_elements(102);
      gj_convolve_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101: marked-successors 
    -- CP-element group 101: 	85 
    -- CP-element group 101: 	89 
    -- CP-element group 101: 	64 
    -- CP-element group 101: 	97 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_update_start_
      -- CP-element group 101: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_Sample/ack
      -- CP-element group 101: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_Update/req
      -- 
    ack_4155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1863_inst_ack_0, ack => convolve_CP_3851_elements(101)); -- 
    req_4159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(101), ack => WPIPE_kernel_pipe1_1863_inst_req_1); -- 
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	140 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	100 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe1_1863_Update/ack
      -- 
    ack_4160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1863_inst_ack_1, ack => convolve_CP_3851_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: 	87 
    -- CP-element group 103: 	91 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	105 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_Sample/req
      -- 
    req_4168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(103), ack => WPIPE_kernel_pipe2_1867_inst_req_0); -- 
    convolve_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(66) & convolve_CP_3851_elements(87) & convolve_CP_3851_elements(91) & convolve_CP_3851_elements(105);
      gj_convolve_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: marked-successors 
    -- CP-element group 104: 	85 
    -- CP-element group 104: 	89 
    -- CP-element group 104: 	64 
    -- CP-element group 104:  members (6) 
      -- CP-element group 104: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_Sample/ack
      -- CP-element group 104: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_Update/req
      -- 
    ack_4169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_1867_inst_ack_0, ack => convolve_CP_3851_elements(104)); -- 
    req_4173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(104), ack => WPIPE_kernel_pipe2_1867_inst_req_1); -- 
    -- CP-element group 105:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	140 
    -- CP-element group 105: marked-successors 
    -- CP-element group 105: 	103 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_kernel_pipe2_1867_Update/ack
      -- 
    ack_4174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_1867_inst_ack_1, ack => convolve_CP_3851_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	66 
    -- CP-element group 106: 	95 
    -- CP-element group 106: 	30 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	108 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_Sample/req
      -- 
    req_4182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(106), ack => WPIPE_input_done_pipe_1888_inst_req_0); -- 
    convolve_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(66) & convolve_CP_3851_elements(95) & convolve_CP_3851_elements(30) & convolve_CP_3851_elements(108);
      gj_convolve_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	26 
    -- CP-element group 107: 	93 
    -- CP-element group 107: 	64 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_update_start_
      -- CP-element group 107: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_Sample/ack
      -- CP-element group 107: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_Update/req
      -- 
    ack_4183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1888_inst_ack_0, ack => convolve_CP_3851_elements(107)); -- 
    req_4187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(107), ack => WPIPE_input_done_pipe_1888_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	140 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	106 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_input_done_pipe_1888_Update/ack
      -- 
    ack_4188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1888_inst_ack_1, ack => convolve_CP_3851_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	49 
    -- CP-element group 109: 	83 
    -- CP-element group 109: 	87 
    -- CP-element group 109: 	91 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_Sample/rr
      -- 
    rr_4196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(109), ack => slice_1893_inst_req_0); -- 
    convolve_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(49) & convolve_CP_3851_elements(83) & convolve_CP_3851_elements(87) & convolve_CP_3851_elements(91) & convolve_CP_3851_elements(111);
      gj_convolve_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	123 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_Update/cr
      -- 
    cr_4201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(110), ack => slice_1893_inst_req_1); -- 
    convolve_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(123) & convolve_CP_3851_elements(112);
      gj_convolve_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	81 
    -- CP-element group 111: 	85 
    -- CP-element group 111: 	89 
    -- CP-element group 111: 	45 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_Sample/ra
      -- 
    ra_4197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1893_inst_ack_0, ack => convolve_CP_3851_elements(111)); -- 
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	121 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1893_Update/ca
      -- 
    ca_4202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1893_inst_ack_1, ack => convolve_CP_3851_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	49 
    -- CP-element group 113: 	83 
    -- CP-element group 113: 	87 
    -- CP-element group 113: 	91 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_Sample/rr
      -- 
    rr_4210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(113), ack => slice_1897_inst_req_0); -- 
    convolve_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(49) & convolve_CP_3851_elements(83) & convolve_CP_3851_elements(87) & convolve_CP_3851_elements(91) & convolve_CP_3851_elements(115);
      gj_convolve_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: 	134 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_update_start_
      -- CP-element group 114: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_Update/cr
      -- 
    cr_4215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(114), ack => slice_1897_inst_req_1); -- 
    convolve_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(116) & convolve_CP_3851_elements(134);
      gj_convolve_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	81 
    -- CP-element group 115: 	85 
    -- CP-element group 115: 	89 
    -- CP-element group 115: 	45 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_Sample/ra
      -- 
    ra_4211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1897_inst_ack_0, ack => convolve_CP_3851_elements(115)); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	132 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/slice_1897_Update/ca
      -- 
    ca_4216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1897_inst_ack_1, ack => convolve_CP_3851_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	95 
    -- CP-element group 117: 	30 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_Sample/req
      -- 
    req_4224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(117), ack => W_next_sum_1872_delayed_1_0_1899_inst_req_0); -- 
    convolve_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(95) & convolve_CP_3851_elements(30) & convolve_CP_3851_elements(119);
      gj_convolve_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: 	123 
    -- CP-element group 118: 	126 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_update_start_
      -- CP-element group 118: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_Update/req
      -- 
    req_4229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(118), ack => W_next_sum_1872_delayed_1_0_1899_inst_req_1); -- 
    convolve_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(120) & convolve_CP_3851_elements(123) & convolve_CP_3851_elements(126);
      gj_convolve_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	26 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	93 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_Sample/ack
      -- 
    ack_4225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1872_delayed_1_0_1899_inst_ack_0, ack => convolve_CP_3851_elements(119)); -- 
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: 	125 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1901_Update/ack
      -- 
    ack_4230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1872_delayed_1_0_1899_inst_ack_1, ack => convolve_CP_3851_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: 	112 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_Sample/rr
      -- 
    rr_4238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(121), ack => type_cast_1905_inst_req_0); -- 
    convolve_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(120) & convolve_CP_3851_elements(112) & convolve_CP_3851_elements(123);
      gj_convolve_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: 	126 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_update_start_
      -- CP-element group 122: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_Update/cr
      -- 
    cr_4243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(122), ack => type_cast_1905_inst_req_1); -- 
    convolve_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(124) & convolve_CP_3851_elements(126);
      gj_convolve_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	110 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_Sample/ra
      -- 
    ra_4239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1905_inst_ack_0, ack => convolve_CP_3851_elements(123)); -- 
    -- CP-element group 124:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124: marked-successors 
    -- CP-element group 124: 	122 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1905_Update/ca
      -- 
    ca_4244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1905_inst_ack_1, ack => convolve_CP_3851_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	120 
    -- CP-element group 125: 	124 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	138 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_Sample/req
      -- 
    req_4252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(125), ack => WPIPE_maxpool_output_pipe_1903_inst_req_0); -- 
    convolve_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(120) & convolve_CP_3851_elements(124) & convolve_CP_3851_elements(138) & convolve_CP_3851_elements(127);
      gj_convolve_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	122 
    -- CP-element group 126: 	118 
    -- CP-element group 126:  members (6) 
      -- CP-element group 126: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_update_start_
      -- CP-element group 126: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_Sample/ack
      -- CP-element group 126: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_Update/req
      -- 
    ack_4253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1903_inst_ack_0, ack => convolve_CP_3851_elements(126)); -- 
    req_4257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(126), ack => WPIPE_maxpool_output_pipe_1903_inst_req_1); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	136 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1903_Update/ack
      -- 
    ack_4258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1903_inst_ack_1, ack => convolve_CP_3851_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	95 
    -- CP-element group 128: 	30 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_Sample/req
      -- 
    req_4266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(128), ack => W_next_sum_1877_delayed_1_0_1907_inst_req_0); -- 
    convolve_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(95) & convolve_CP_3851_elements(30) & convolve_CP_3851_elements(130);
      gj_convolve_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	137 
    -- CP-element group 129: 	131 
    -- CP-element group 129: 	134 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_update_start_
      -- CP-element group 129: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_Update/req
      -- 
    req_4271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(129), ack => W_next_sum_1877_delayed_1_0_1907_inst_req_1); -- 
    convolve_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(137) & convolve_CP_3851_elements(131) & convolve_CP_3851_elements(134);
      gj_convolve_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	26 
    -- CP-element group 130: 	128 
    -- CP-element group 130: 	93 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_Sample/ack
      -- 
    ack_4267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1877_delayed_1_0_1907_inst_ack_0, ack => convolve_CP_3851_elements(130)); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	136 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/assign_stmt_1909_Update/ack
      -- 
    ack_4272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1877_delayed_1_0_1907_inst_ack_1, ack => convolve_CP_3851_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	116 
    -- CP-element group 132: 	131 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_Sample/rr
      -- 
    rr_4280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(132), ack => type_cast_1913_inst_req_0); -- 
    convolve_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(116) & convolve_CP_3851_elements(131) & convolve_CP_3851_elements(134);
      gj_convolve_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	137 
    -- CP-element group 133: 	135 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_update_start_
      -- CP-element group 133: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_Update/cr
      -- 
    cr_4285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(133), ack => type_cast_1913_inst_req_1); -- 
    convolve_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(137) & convolve_CP_3851_elements(135);
      gj_convolve_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	114 
    -- CP-element group 134: 	129 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_Sample/ra
      -- 
    ra_4281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1913_inst_ack_0, ack => convolve_CP_3851_elements(134)); -- 
    -- CP-element group 135:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/type_cast_1913_Update/ca
      -- 
    ca_4286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1913_inst_ack_1, ack => convolve_CP_3851_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	127 
    -- CP-element group 136: 	131 
    -- CP-element group 136: 	135 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_Sample/req
      -- 
    req_4294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(136), ack => WPIPE_maxpool_output_pipe_1911_inst_req_0); -- 
    convolve_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(127) & convolve_CP_3851_elements(131) & convolve_CP_3851_elements(135) & convolve_CP_3851_elements(138);
      gj_convolve_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	129 
    -- CP-element group 137: 	133 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_update_start_
      -- CP-element group 137: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_Sample/ack
      -- CP-element group 137: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_Update/req
      -- 
    ack_4295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1911_inst_ack_0, ack => convolve_CP_3851_elements(137)); -- 
    req_4299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(137), ack => WPIPE_maxpool_output_pipe_1911_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	125 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/WPIPE_maxpool_output_pipe_1911_Update/ack
      -- 
    ack_4300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1911_inst_ack_1, ack => convolve_CP_3851_elements(138)); -- 
    -- CP-element group 139:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	19 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	20 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_3851_elements(139) is a control-delay.
    cp_element_139_delay: control_delay_element  generic map(name => " 139_delay", delay_value => 1)  port map(req => convolve_CP_3851_elements(19), ack => convolve_CP_3851_elements(139), clk => clk, reset =>reset);
    -- CP-element group 140:  join  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: 	102 
    -- CP-element group 140: 	105 
    -- CP-element group 140: 	108 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	16 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_1739/do_while_stmt_1764/do_while_stmt_1764_loop_body/$exit
      -- 
    convolve_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_3851_elements(138) & convolve_CP_3851_elements(102) & convolve_CP_3851_elements(105) & convolve_CP_3851_elements(108);
      gj_convolve_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_3851_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	15 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_1739/do_while_stmt_1764/loop_exit/$exit
      -- CP-element group 141: 	 branch_block_stmt_1739/do_while_stmt_1764/loop_exit/ack
      -- 
    ack_4305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1764_branch_ack_0, ack => convolve_CP_3851_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	15 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1739/do_while_stmt_1764/loop_taken/$exit
      -- CP-element group 142: 	 branch_block_stmt_1739/do_while_stmt_1764/loop_taken/ack
      -- 
    ack_4309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1764_branch_ack_1, ack => convolve_CP_3851_elements(142)); -- 
    -- CP-element group 143:  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	13 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	2 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1739/do_while_stmt_1764/$exit
      -- 
    convolve_CP_3851_elements(143) <= convolve_CP_3851_elements(13);
    -- CP-element group 144:  merge  fork  transition  place  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	0 
    -- CP-element group 144: 	2 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	10 
    -- CP-element group 144: 	3 
    -- CP-element group 144: 	5 
    -- CP-element group 144: 	8 
    -- CP-element group 144:  members (19) 
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_Update/cr
      -- CP-element group 144: 	 branch_block_stmt_1739/merge_stmt_1740__exit__
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763__entry__
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/$entry
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_num_out_pipe_1742_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/RPIPE_size_pipe_1745_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_update_start_
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1749_Update/cr
      -- CP-element group 144: 	 branch_block_stmt_1739/assign_stmt_1743_to_assign_stmt_1763/slice_1753_update_start_
      -- CP-element group 144: 	 branch_block_stmt_1739/merge_stmt_1740_PhiReqMerge
      -- CP-element group 144: 	 branch_block_stmt_1739/merge_stmt_1740_PhiAck/$entry
      -- CP-element group 144: 	 branch_block_stmt_1739/merge_stmt_1740_PhiAck/$exit
      -- CP-element group 144: 	 branch_block_stmt_1739/merge_stmt_1740_PhiAck/dummy
      -- 
    cr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(144), ack => slice_1753_inst_req_1); -- 
    rr_3876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(144), ack => RPIPE_num_out_pipe_1742_inst_req_0); -- 
    rr_3890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(144), ack => RPIPE_size_pipe_1745_inst_req_0); -- 
    cr_3909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_3851_elements(144), ack => slice_1749_inst_req_1); -- 
    convolve_CP_3851_elements(144) <= OrReduce(convolve_CP_3851_elements(0) & convolve_CP_3851_elements(2));
    convolve_do_while_stmt_1764_terminator_4310: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_1764_terminator_4310", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_3851_elements(16),loop_continue => convolve_CP_3851_elements(142),loop_terminate => convolve_CP_3851_elements(141),loop_back => convolve_CP_3851_elements(14),loop_exit => convolve_CP_3851_elements(13),clk => clk, reset => reset); -- 
    phi_stmt_1766_phi_seq_3988_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3851_elements(31);
      convolve_CP_3851_elements(36)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3851_elements(38);
      convolve_CP_3851_elements(37)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3851_elements(39);
      convolve_CP_3851_elements(32) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3851_elements(33);
      convolve_CP_3851_elements(40)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3851_elements(40);
      convolve_CP_3851_elements(41)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3851_elements(42);
      convolve_CP_3851_elements(34) <= phi_mux_reqs(1);
      phi_stmt_1766_phi_seq_3988 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1766_phi_seq_3988") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3851_elements(27), 
          phi_sample_ack => convolve_CP_3851_elements(28), 
          phi_update_req => convolve_CP_3851_elements(29), 
          phi_update_ack => convolve_CP_3851_elements(30), 
          phi_mux_ack => convolve_CP_3851_elements(35), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1770_phi_seq_4032_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3851_elements(50);
      convolve_CP_3851_elements(55)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3851_elements(57);
      convolve_CP_3851_elements(56)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3851_elements(58);
      convolve_CP_3851_elements(51) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3851_elements(52);
      convolve_CP_3851_elements(59)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3851_elements(59);
      convolve_CP_3851_elements(60)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3851_elements(61);
      convolve_CP_3851_elements(53) <= phi_mux_reqs(1);
      phi_stmt_1770_phi_seq_4032 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1770_phi_seq_4032") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3851_elements(46), 
          phi_sample_ack => convolve_CP_3851_elements(47), 
          phi_update_req => convolve_CP_3851_elements(48), 
          phi_update_ack => convolve_CP_3851_elements(49), 
          phi_mux_ack => convolve_CP_3851_elements(54), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1774_phi_seq_4076_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_3851_elements(69);
      convolve_CP_3851_elements(72)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_3851_elements(72);
      convolve_CP_3851_elements(73)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_3851_elements(74);
      convolve_CP_3851_elements(70) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_3851_elements(67);
      convolve_CP_3851_elements(76)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_3851_elements(78);
      convolve_CP_3851_elements(77)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_3851_elements(79);
      convolve_CP_3851_elements(68) <= phi_mux_reqs(1);
      phi_stmt_1774_phi_seq_4076 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1774_phi_seq_4076") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_3851_elements(21), 
          phi_sample_ack => convolve_CP_3851_elements(65), 
          phi_update_req => convolve_CP_3851_elements(23), 
          phi_update_ack => convolve_CP_3851_elements(66), 
          phi_mux_ack => convolve_CP_3851_elements(71), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3940_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_3851_elements(17);
        preds(1)  <= convolve_CP_3851_elements(18);
        entry_tmerge_3940 : transition_merge -- 
          generic map(name => " entry_tmerge_3940")
          port map (preds => preds, symbol_out => convolve_CP_3851_elements(19));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_1877_wire : std_logic_vector(15 downto 0);
    signal ADD_u31_u31_1838_wire : std_logic_vector(30 downto 0);
    signal MUX_1878_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_1826_1826_delayed_1_0_1849 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1852_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1858_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1917_wire : std_logic_vector(0 downto 0);
    signal SUB_u31_u31_1793_1793_delayed_1_0_1814 : std_logic_vector(30 downto 0);
    signal acc_1770 : std_logic_vector(15 downto 0);
    signal acc_val_1826 : std_logic_vector(15 downto 0);
    signal acc_val_dn_1898 : std_logic_vector(7 downto 0);
    signal acc_val_up_1894 : std_logic_vector(7 downto 0);
    signal acc_var_1763 : std_logic_vector(15 downto 0);
    signal all_done_flag_1886 : std_logic_vector(0 downto 0);
    signal iread_1782 : std_logic_vector(15 downto 0);
    signal ival_1786 : std_logic_vector(15 downto 0);
    signal konst_1812_wire_constant : std_logic_vector(30 downto 0);
    signal konst_1829_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1835_wire_constant : std_logic_vector(30 downto 0);
    signal konst_1837_wire_constant : std_logic_vector(30 downto 0);
    signal konst_1876_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1889_wire_constant : std_logic_vector(0 downto 0);
    signal kread_1800 : std_logic_vector(15 downto 0);
    signal kval_1804 : std_logic_vector(15 downto 0);
    signal mcount_var_1758 : std_logic_vector(30 downto 0);
    signal mul_val_1809 : std_logic_vector(15 downto 0);
    signal mycount_1766 : std_logic_vector(30 downto 0);
    signal n_out_count_1881 : std_logic_vector(15 downto 0);
    signal n_out_count_1881_1778_buffered : std_logic_vector(15 downto 0);
    signal nacc_1832 : std_logic_vector(15 downto 0);
    signal nacc_1832_1772_buffered : std_logic_vector(15 downto 0);
    signal next_sum_1819 : std_logic_vector(0 downto 0);
    signal next_sum_1872_delayed_1_0_1901 : std_logic_vector(0 downto 0);
    signal next_sum_1877_delayed_1_0_1909 : std_logic_vector(0 downto 0);
    signal nmycount_1840 : std_logic_vector(30 downto 0);
    signal nmycount_1840_1768_buffered : std_logic_vector(30 downto 0);
    signal num_out_1743 : std_logic_vector(15 downto 0);
    signal out_count_1774 : std_logic_vector(15 downto 0);
    signal out_done_flag_1845 : std_logic_vector(0 downto 0);
    signal pingpong_1750 : std_logic_vector(0 downto 0);
    signal send_back1_1855 : std_logic_vector(0 downto 0);
    signal send_back2_1861 : std_logic_vector(0 downto 0);
    signal size_1754 : std_logic_vector(30 downto 0);
    signal size_read_1746 : std_logic_vector(31 downto 0);
    signal temp1_1790 : std_logic_vector(15 downto 0);
    signal temp2_1794 : std_logic_vector(15 downto 0);
    signal type_cast_1777_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1822_wire : std_logic_vector(15 downto 0);
    signal type_cast_1824_wire : std_logic_vector(15 downto 0);
    signal type_cast_1874_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1905_wire : std_logic_vector(7 downto 0);
    signal type_cast_1913_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    acc_var_1763 <= "0000000000000000";
    konst_1812_wire_constant <= "0000000000000000000000000000001";
    konst_1829_wire_constant <= "0000000000000000";
    konst_1835_wire_constant <= "0000000000000000000000000000000";
    konst_1837_wire_constant <= "0000000000000000000000000000001";
    konst_1876_wire_constant <= "0000000000000001";
    konst_1889_wire_constant <= "1";
    mcount_var_1758 <= "0000000000000000000000000000000";
    type_cast_1777_wire_constant <= "0000000000000001";
    type_cast_1874_wire_constant <= "0000000000000001";
    phi_stmt_1766: Block -- phi operator 
      signal idata: std_logic_vector(61 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_1840_1768_buffered & mcount_var_1758;
      req <= phi_stmt_1766_req_0 & phi_stmt_1766_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1766",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 31) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1766_ack_0,
          idata => idata,
          odata => mycount_1766,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1766
    phi_stmt_1770: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nacc_1832_1772_buffered & acc_var_1763;
      req <= phi_stmt_1770_req_0 & phi_stmt_1770_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1770",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1770_ack_0,
          idata => idata,
          odata => acc_1770,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1770
    phi_stmt_1774: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1777_wire_constant & n_out_count_1881_1778_buffered;
      req <= phi_stmt_1774_req_0 & phi_stmt_1774_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1774",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1774_ack_0,
          idata => idata,
          odata => out_count_1774,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1774
    -- flow-through select operator MUX_1799_inst
    kread_1800 <= temp2_1794 when (pingpong_1750(0) /=  '0') else temp1_1790;
    -- flow-through select operator MUX_1831_inst
    nacc_1832 <= konst_1829_wire_constant when (next_sum_1819(0) /=  '0') else acc_val_1826;
    -- flow-through select operator MUX_1839_inst
    nmycount_1840 <= konst_1835_wire_constant when (next_sum_1819(0) /=  '0') else ADD_u31_u31_1838_wire;
    -- flow-through select operator MUX_1878_inst
    MUX_1878_wire <= type_cast_1874_wire_constant when (out_done_flag_1845(0) /=  '0') else ADD_u16_u16_1877_wire;
    -- flow-through select operator MUX_1880_inst
    n_out_count_1881 <= MUX_1878_wire when (next_sum_1819(0) /=  '0') else out_count_1774;
    slice_1749_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1749_inst_req_0;
      slice_1749_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1749_inst_req_1;
      slice_1749_inst_ack_1<= update_ack(0);
      slice_1749_inst: SliceSplitProtocol generic map(name => "slice_1749_inst", in_data_width => 32, high_index => 31, low_index => 31, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => size_read_1746, dout => pingpong_1750, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1753_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1753_inst_req_0;
      slice_1753_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1753_inst_req_1;
      slice_1753_inst_ack_1<= update_ack(0);
      slice_1753_inst: SliceSplitProtocol generic map(name => "slice_1753_inst", in_data_width => 32, high_index => 30, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => size_read_1746, dout => size_1754, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1893_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1893_inst_req_0;
      slice_1893_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1893_inst_req_1;
      slice_1893_inst_ack_1<= update_ack(0);
      slice_1893_inst: SliceSplitProtocol generic map(name => "slice_1893_inst", in_data_width => 16, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1826, dout => acc_val_up_1894, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1897_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1897_inst_req_0;
      slice_1897_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1897_inst_req_1;
      slice_1897_inst_ack_1<= update_ack(0);
      slice_1897_inst: SliceSplitProtocol generic map(name => "slice_1897_inst", in_data_width => 16, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1826, dout => acc_val_dn_1898, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_next_sum_1872_delayed_1_0_1899_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1872_delayed_1_0_1899_inst_req_0;
      W_next_sum_1872_delayed_1_0_1899_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1872_delayed_1_0_1899_inst_req_1;
      W_next_sum_1872_delayed_1_0_1899_inst_ack_1<= rack(0);
      W_next_sum_1872_delayed_1_0_1899_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1872_delayed_1_0_1899_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1872_delayed_1_0_1901,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_next_sum_1877_delayed_1_0_1907_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1877_delayed_1_0_1907_inst_req_0;
      W_next_sum_1877_delayed_1_0_1907_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1877_delayed_1_0_1907_inst_req_1;
      W_next_sum_1877_delayed_1_0_1907_inst_ack_1<= rack(0);
      W_next_sum_1877_delayed_1_0_1907_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1877_delayed_1_0_1907_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1877_delayed_1_0_1909,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_out_count_1881_1778_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_out_count_1881_1778_buf_req_0;
      n_out_count_1881_1778_buf_ack_0<= wack(0);
      rreq(0) <= n_out_count_1881_1778_buf_req_1;
      n_out_count_1881_1778_buf_ack_1<= rack(0);
      n_out_count_1881_1778_buf : InterlockBuffer generic map ( -- 
        name => "n_out_count_1881_1778_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_out_count_1881,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_out_count_1881_1778_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc_1832_1772_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc_1832_1772_buf_req_0;
      nacc_1832_1772_buf_ack_0<= wack(0);
      rreq(0) <= nacc_1832_1772_buf_req_1;
      nacc_1832_1772_buf_ack_1<= rack(0);
      nacc_1832_1772_buf : InterlockBuffer generic map ( -- 
        name => "nacc_1832_1772_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc_1832,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc_1832_1772_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_1840_1768_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_1840_1768_buf_req_0;
      nmycount_1840_1768_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_1840_1768_buf_req_1;
      nmycount_1840_1768_buf_ack_1<= rack(0);
      nmycount_1840_1768_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_1840_1768_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 31,
        out_data_width => 31,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_1840,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_1840_1768_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1785_inst
    process(iread_1782) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread_1782(15 downto 0);
      ival_1786 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1803_inst
    process(kread_1800) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread_1800(15 downto 0);
      kval_1804 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1822_inst
    process(acc_1770) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := acc_1770(15 downto 0);
      type_cast_1822_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1824_inst
    process(mul_val_1809) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := mul_val_1809(15 downto 0);
      type_cast_1824_wire <= tmp_var; -- 
    end process;
    type_cast_1905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1905_inst_req_0;
      type_cast_1905_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1905_inst_req_1;
      type_cast_1905_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1872_delayed_1_0_1901(0);
      type_cast_1905_inst_gI: SplitGuardInterface generic map(name => "type_cast_1905_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1905_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1905_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_up_1894,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1905_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1913_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1913_inst_req_0;
      type_cast_1913_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1913_inst_req_1;
      type_cast_1913_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1877_delayed_1_0_1909(0);
      type_cast_1913_inst_gI: SplitGuardInterface generic map(name => "type_cast_1913_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1913_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1913_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_dn_1898,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1913_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1764_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1917_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1764_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1764_branch_req_0,
          ack0 => do_while_stmt_1764_branch_ack_0,
          ack1 => do_while_stmt_1764_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_1825_inst
    process(type_cast_1822_wire, type_cast_1824_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_1822_wire, type_cast_1824_wire, tmp_var);
      acc_val_1826 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1877_inst
    process(out_count_1774) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(out_count_1774, konst_1876_wire_constant, tmp_var);
      ADD_u16_u16_1877_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u31_u31_1838_inst
    process(mycount_1766) -- 
      variable tmp_var : std_logic_vector(30 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_1766, konst_1837_wire_constant, tmp_var);
      ADD_u31_u31_1838_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1854_inst
    process(NOT_u1_u1_1852_wire, NOT_u1_u1_1826_1826_delayed_1_0_1849) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1852_wire, NOT_u1_u1_1826_1826_delayed_1_0_1849, tmp_var);
      send_back1_1855 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1860_inst
    process(NOT_u1_u1_1858_wire, pingpong_1750) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1858_wire, pingpong_1750, tmp_var);
      send_back2_1861 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1885_inst
    process(out_done_flag_1845, next_sum_1819) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_1845, next_sum_1819, tmp_var);
      all_done_flag_1886 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1844_inst
    process(out_count_1774, num_out_1743) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(out_count_1774, num_out_1743, tmp_var);
      out_done_flag_1845 <= tmp_var; --
    end process;
    -- binary operator EQ_u31_u1_1818_inst
    process(mycount_1766, SUB_u31_u31_1793_1793_delayed_1_0_1814) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycount_1766, SUB_u31_u31_1793_1793_delayed_1_0_1814, tmp_var);
      next_sum_1819 <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_1808_inst
    process(kval_1804, ival_1786) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval_1804, ival_1786, tmp_var);
      mul_val_1809 <= tmp_var; --
    end process;
    -- shared split operator group (9) : NOT_u1_u1_1848_inst 
    ApIntNot_group_9: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pingpong_1750;
      NOT_u1_u1_1826_1826_delayed_1_0_1849 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1848_inst_req_0;
      NOT_u1_u1_1848_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1848_inst_req_1;
      NOT_u1_u1_1848_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_9_gI: SplitGuardInterface generic map(name => "ApIntNot_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- unary operator NOT_u1_u1_1852_inst
    process(out_done_flag_1845) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", out_done_flag_1845, tmp_var);
      NOT_u1_u1_1852_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1858_inst
    process(out_done_flag_1845) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", out_done_flag_1845, tmp_var);
      NOT_u1_u1_1858_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1917_inst
    process(all_done_flag_1886) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", all_done_flag_1886, tmp_var);
      NOT_u1_u1_1917_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (13) : SUB_u31_u31_1813_inst 
    ApIntSub_group_13: Block -- 
      signal data_in: std_logic_vector(30 downto 0);
      signal data_out: std_logic_vector(30 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= size_1754;
      SUB_u31_u31_1793_1793_delayed_1_0_1814 <= data_out(30 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u31_u31_1813_inst_req_0;
      SUB_u31_u31_1813_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u31_u31_1813_inst_req_1;
      SUB_u31_u31_1813_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_13_gI: SplitGuardInterface generic map(name => "ApIntSub_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 31,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 31,
          constant_operand => "0000000000000000000000000000001",
          constant_width => 31,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared inport operator group (0) : RPIPE_input_pipe1_1781_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_1781_inst_req_0;
      RPIPE_input_pipe1_1781_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_1781_inst_req_1;
      RPIPE_input_pipe1_1781_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iread_1782 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_kernel_pipe1_1789_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_1789_inst_req_0;
      RPIPE_kernel_pipe1_1789_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_1789_inst_req_1;
      RPIPE_kernel_pipe1_1789_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not pingpong_1750(0);
      temp1_1790 <= data_out(15 downto 0);
      kernel_pipe1_read_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_1: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_kernel_pipe2_1793_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe2_1793_inst_req_0;
      RPIPE_kernel_pipe2_1793_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe2_1793_inst_req_1;
      RPIPE_kernel_pipe2_1793_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= pingpong_1750(0);
      temp2_1794 <= data_out(15 downto 0);
      kernel_pipe2_read_2_gI: SplitGuardInterface generic map(name => "kernel_pipe2_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_read_2: InputPortRevised -- 
        generic map ( name => "kernel_pipe2_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe2_pipe_read_req(0),
          oack => kernel_pipe2_pipe_read_ack(0),
          odata => kernel_pipe2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_num_out_pipe_1742_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_num_out_pipe_1742_inst_req_0;
      RPIPE_num_out_pipe_1742_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_num_out_pipe_1742_inst_req_1;
      RPIPE_num_out_pipe_1742_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      num_out_1743 <= data_out(15 downto 0);
      num_out_pipe_read_3_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_3: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_size_pipe_1745_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_1745_inst_req_0;
      RPIPE_size_pipe_1745_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_1745_inst_req_1;
      RPIPE_size_pipe_1745_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      size_read_1746 <= data_out(31 downto 0);
      size_pipe_read_4_gI: SplitGuardInterface generic map(name => "size_pipe_read_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_4: InputPortRevised -- 
        generic map ( name => "size_pipe_read_4", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_input_done_pipe_1888_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_1888_inst_req_0;
      WPIPE_input_done_pipe_1888_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_1888_inst_req_1;
      WPIPE_input_done_pipe_1888_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= all_done_flag_1886(0);
      data_in <= konst_1889_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe1_1863_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_1863_inst_req_0;
      WPIPE_kernel_pipe1_1863_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_1863_inst_req_1;
      WPIPE_kernel_pipe1_1863_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_back1_1855(0);
      data_in <= kread_1800;
      kernel_pipe1_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_kernel_pipe2_1867_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe2_1867_inst_req_0;
      WPIPE_kernel_pipe2_1867_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe2_1867_inst_req_1;
      WPIPE_kernel_pipe2_1867_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_back2_1861(0);
      data_in <= kread_1800;
      kernel_pipe2_write_2_gI: SplitGuardInterface generic map(name => "kernel_pipe2_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_write_2: OutputPortRevised -- 
        generic map ( name => "kernel_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe2_pipe_write_req(0),
          oack => kernel_pipe2_pipe_write_ack(0),
          odata => kernel_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_maxpool_output_pipe_1911_inst WPIPE_maxpool_output_pipe_1903_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1911_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1903_inst_req_0;
      WPIPE_maxpool_output_pipe_1911_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1903_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1911_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1903_inst_req_1;
      WPIPE_maxpool_output_pipe_1911_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1903_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= next_sum_1872_delayed_1_0_1901(0);
      guard_vector(1)  <= next_sum_1877_delayed_1_0_1909(0);
      data_in <= type_cast_1913_wire & type_cast_1905_wire;
      maxpool_output_pipe_write_3_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_3: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    end_add : in  std_logic_vector(63 downto 0);
    pp : in  std_logic_vector(7 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 136)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal end_add_buffer :  std_logic_vector(63 downto 0);
  signal end_add_update_enable: Boolean;
  signal pp_buffer :  std_logic_vector(7 downto 0);
  signal pp_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_671_start: Boolean;
  signal loadKernelChannel_CP_671_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_413_index_offset_ack_0 : boolean;
  signal array_obj_ref_413_index_offset_req_1 : boolean;
  signal do_while_stmt_361_branch_ack_0 : boolean;
  signal W_fetch_val_412_delayed_13_0_427_inst_ack_0 : boolean;
  signal WPIPE_size_pipe_443_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_397_inst_ack_1 : boolean;
  signal W_fn_410_delayed_13_0_424_inst_ack_0 : boolean;
  signal CONCAT_u1_u32_450_inst_req_1 : boolean;
  signal array_obj_ref_413_index_offset_ack_1 : boolean;
  signal WPIPE_size_pipe_443_inst_ack_0 : boolean;
  signal CONCAT_u1_u32_450_inst_ack_0 : boolean;
  signal W_fn_410_delayed_13_0_424_inst_ack_1 : boolean;
  signal CONCAT_u1_u32_450_inst_ack_1 : boolean;
  signal CONCAT_u1_u32_450_inst_req_0 : boolean;
  signal ptr_deref_422_load_0_ack_0 : boolean;
  signal addr_of_414_final_reg_req_0 : boolean;
  signal phi_stmt_367_ack_0 : boolean;
  signal phi_stmt_367_req_0 : boolean;
  signal WPIPE_size_pipe_443_inst_req_1 : boolean;
  signal WPIPE_size_pipe_443_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe2_397_inst_req_1 : boolean;
  signal ptr_deref_422_load_0_req_0 : boolean;
  signal nfetch_val_435_370_buf_ack_1 : boolean;
  signal nfetch_val_435_370_buf_req_1 : boolean;
  signal addr_of_414_final_reg_ack_0 : boolean;
  signal my_fetch_350_369_buf_req_0 : boolean;
  signal phi_stmt_367_req_1 : boolean;
  signal W_fn_410_delayed_13_0_424_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_393_inst_req_0 : boolean;
  signal array_obj_ref_413_index_offset_req_0 : boolean;
  signal addr_of_414_final_reg_req_1 : boolean;
  signal WPIPE_kernel_pipe2_397_inst_ack_0 : boolean;
  signal W_fetch_val_412_delayed_13_0_427_inst_req_1 : boolean;
  signal my_fetch_350_369_buf_ack_0 : boolean;
  signal addr_of_414_final_reg_ack_1 : boolean;
  signal nfetch_val_435_370_buf_req_0 : boolean;
  signal W_fetch_val_412_delayed_13_0_427_inst_ack_1 : boolean;
  signal my_fetch_350_369_buf_req_1 : boolean;
  signal nfetch_val_435_370_buf_ack_0 : boolean;
  signal W_fn_410_delayed_13_0_424_inst_req_1 : boolean;
  signal W_fn_404_delayed_7_0_416_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_393_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_397_inst_req_0 : boolean;
  signal W_fn_404_delayed_7_0_416_inst_ack_0 : boolean;
  signal W_fetch_val_412_delayed_13_0_427_inst_req_0 : boolean;
  signal ptr_deref_422_load_0_req_1 : boolean;
  signal do_while_stmt_361_branch_ack_1 : boolean;
  signal my_fetch_350_369_buf_ack_1 : boolean;
  signal ptr_deref_422_load_0_ack_1 : boolean;
  signal start_add_366_buf_ack_1 : boolean;
  signal array_obj_ref_344_index_offset_req_0 : boolean;
  signal array_obj_ref_344_index_offset_ack_0 : boolean;
  signal array_obj_ref_344_index_offset_req_1 : boolean;
  signal array_obj_ref_344_index_offset_ack_1 : boolean;
  signal addr_of_345_final_reg_req_0 : boolean;
  signal addr_of_345_final_reg_ack_0 : boolean;
  signal addr_of_345_final_reg_req_1 : boolean;
  signal addr_of_345_final_reg_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_393_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_393_inst_req_1 : boolean;
  signal start_add_366_buf_req_1 : boolean;
  signal W_fn_404_delayed_7_0_416_inst_ack_1 : boolean;
  signal W_fn_404_delayed_7_0_416_inst_req_1 : boolean;
  signal ptr_deref_349_load_0_req_0 : boolean;
  signal ptr_deref_349_load_0_ack_0 : boolean;
  signal ptr_deref_349_load_0_req_1 : boolean;
  signal ptr_deref_349_load_0_ack_1 : boolean;
  signal RPIPE_input_done_pipe_358_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_358_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_358_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_358_inst_ack_1 : boolean;
  signal do_while_stmt_361_branch_req_0 : boolean;
  signal phi_stmt_363_req_0 : boolean;
  signal phi_stmt_363_req_1 : boolean;
  signal phi_stmt_363_ack_0 : boolean;
  signal nmycount_385_365_buf_req_0 : boolean;
  signal nmycount_385_365_buf_ack_0 : boolean;
  signal nmycount_385_365_buf_req_1 : boolean;
  signal nmycount_385_365_buf_ack_1 : boolean;
  signal start_add_366_buf_req_0 : boolean;
  signal start_add_366_buf_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 136) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(127 downto 64) <= end_add;
  end_add_buffer <= in_buffer_data_out(127 downto 64);
  in_buffer_data_in(135 downto 128) <= pp;
  pp_buffer <= in_buffer_data_out(135 downto 128);
  in_buffer_data_in(tag_length + 135 downto 136) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 135 downto 136);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_671_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_671_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_671_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_671_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_671: Block -- control-path 
    signal loadKernelChannel_CP_671_elements: BooleanArray(97 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_671_elements(0) <= loadKernelChannel_CP_671_start;
    loadKernelChannel_CP_671_symbol <= loadKernelChannel_CP_671_elements(97);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/$entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_update_start_
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_resized_1
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_computed_1
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_complete/$entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_complete/req
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_update_start_
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/$entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_sample_start_
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_Sample/rr
      -- 
    cr_766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => ptr_deref_349_load_0_req_1); -- 
    req_701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => array_obj_ref_344_index_offset_req_0); -- 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => array_obj_ref_344_index_offset_req_1); -- 
    rr_780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => RPIPE_input_done_pipe_358_inst_req_0); -- 
    req_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => addr_of_345_final_reg_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_final_index_sum_regn_Sample/ack
      -- 
    ack_702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_344_index_offset_ack_0, ack => loadKernelChannel_CP_671_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_sample_start_
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_offset_calculated
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/array_obj_ref_344_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_request/$entry
      -- CP-element group 2: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_request/req
      -- 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_344_index_offset_ack_1, ack => loadKernelChannel_CP_671_elements(2)); -- 
    req_716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(2), ack => addr_of_345_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_sample_completed_
      -- CP-element group 3: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_request/$exit
      -- CP-element group 3: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_request/ack
      -- 
    ack_717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_345_final_reg_ack_0, ack => loadKernelChannel_CP_671_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_update_completed_
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_complete/$exit
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/addr_of_345_complete/ack
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_sample_start_
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_base_address_resized
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Sample/word_access_start/word_0/rr
      -- 
    ack_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_345_final_reg_ack_1, ack => loadKernelChannel_CP_671_elements(4)); -- 
    rr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(4), ack => ptr_deref_349_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_sample_completed_
      -- CP-element group 5: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Sample/word_access_start/word_0/ra
      -- 
    ra_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_349_load_0_ack_0, ack => loadKernelChannel_CP_671_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_update_completed_
      -- CP-element group 6: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/$exit
      -- CP-element group 6: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/ptr_deref_349_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/ptr_deref_349_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/ptr_deref_349_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_335_to_assign_stmt_359/ptr_deref_349_Update/ptr_deref_349_Merge/merge_ack
      -- 
    ca_767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_349_load_0_ack_1, ack => loadKernelChannel_CP_671_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_sample_completed_
      -- CP-element group 7: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_update_start_
      -- CP-element group 7: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_Sample/ra
      -- CP-element group 7: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_Update/$entry
      -- CP-element group 7: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_Update/cr
      -- 
    ra_781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_358_inst_ack_0, ack => loadKernelChannel_CP_671_elements(7)); -- 
    cr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(7), ack => RPIPE_input_done_pipe_358_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_update_completed_
      -- CP-element group 8: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_Update/$exit
      -- CP-element group 8: 	 assign_stmt_335_to_assign_stmt_359/RPIPE_input_done_pipe_358_Update/ca
      -- 
    ca_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_358_inst_ack_1, ack => loadKernelChannel_CP_671_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	8 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 assign_stmt_335_to_assign_stmt_359/$exit
      -- CP-element group 9: 	 branch_block_stmt_360/$entry
      -- CP-element group 9: 	 branch_block_stmt_360/branch_block_stmt_360__entry__
      -- CP-element group 9: 	 branch_block_stmt_360/do_while_stmt_361__entry__
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(1) & loadKernelChannel_CP_671_elements(8) & loadKernelChannel_CP_671_elements(6);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	93 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	94 
    -- CP-element group 10: 	95 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 assign_stmt_451/CONCAT_u1_u32_450_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_451/CONCAT_u1_u32_450_Update/cr
      -- CP-element group 10: 	 assign_stmt_451/CONCAT_u1_u32_450_Sample/rr
      -- CP-element group 10: 	 assign_stmt_451/CONCAT_u1_u32_450_Update/$entry
      -- CP-element group 10: 	 assign_stmt_451/CONCAT_u1_u32_450_sample_start_
      -- CP-element group 10: 	 assign_stmt_451/$entry
      -- CP-element group 10: 	 assign_stmt_451/CONCAT_u1_u32_450_update_start_
      -- CP-element group 10: 	 branch_block_stmt_360/$exit
      -- CP-element group 10: 	 branch_block_stmt_360/branch_block_stmt_360__exit__
      -- CP-element group 10: 	 branch_block_stmt_360/do_while_stmt_361__exit__
      -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(10), ack => CONCAT_u1_u32_450_inst_req_1); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(10), ack => CONCAT_u1_u32_450_inst_req_0); -- 
    loadKernelChannel_CP_671_elements(10) <= loadKernelChannel_CP_671_elements(93);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_360/do_while_stmt_361/$entry
      -- CP-element group 11: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361__entry__
      -- 
    loadKernelChannel_CP_671_elements(11) <= loadKernelChannel_CP_671_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	93 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361__exit__
      -- 
    -- Element group loadKernelChannel_CP_671_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_360/do_while_stmt_361/loop_back
      -- 
    -- Element group loadKernelChannel_CP_671_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	91 
    -- CP-element group 14: 	92 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_360/do_while_stmt_361/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_360/do_while_stmt_361/loop_taken/$entry
      -- CP-element group 14: 	 branch_block_stmt_360/do_while_stmt_361/condition_done
      -- 
    loadKernelChannel_CP_671_elements(14) <= loadKernelChannel_CP_671_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	90 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_360/do_while_stmt_361/loop_body_done
      -- 
    loadKernelChannel_CP_671_elements(15) <= loadKernelChannel_CP_671_elements(90);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	47 
    -- CP-element group 16: 	30 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_671_elements(16) <= loadKernelChannel_CP_671_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	49 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_671_elements(17) <= loadKernelChannel_CP_671_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	89 
    -- CP-element group 18: 	67 
    -- CP-element group 18: 	43 
    -- CP-element group 18: 	44 
    -- CP-element group 18: 	68 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	25 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_671_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	89 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	29 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/condition_evaluated
      -- 
    condition_evaluated_808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(19), ack => do_while_stmt_361_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(89) & loadKernelChannel_CP_671_elements(23) & loadKernelChannel_CP_671_elements(29);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	24 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	26 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_sample_start__ps
      -- CP-element group 20: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/aggregated_phi_sample_req
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(43) & loadKernelChannel_CP_671_elements(24) & loadKernelChannel_CP_671_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	45 
    -- CP-element group 21: 	27 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	82 
    -- CP-element group 21: 	78 
    -- CP-element group 21: 	86 
    -- CP-element group 21: 	90 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	43 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(45) & loadKernelChannel_CP_671_elements(27);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	44 
    -- CP-element group 22: 	25 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	28 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/aggregated_phi_update_req
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(44) & loadKernelChannel_CP_671_elements(25);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	46 
    -- CP-element group 23: 	29 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(29);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	75 
    -- CP-element group 25: 	83 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	64 
    -- CP-element group 25: 	69 
    -- CP-element group 25: 	29 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(75) & loadKernelChannel_CP_671_elements(83) & loadKernelChannel_CP_671_elements(61) & loadKernelChannel_CP_671_elements(64) & loadKernelChannel_CP_671_elements(69) & loadKernelChannel_CP_671_elements(29);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	20 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_sample_start__ps
      -- 
    loadKernelChannel_CP_671_elements(26) <= loadKernelChannel_CP_671_elements(20);
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	21 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_671_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	22 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_update_start__ps
      -- 
    loadKernelChannel_CP_671_elements(28) <= loadKernelChannel_CP_671_elements(22);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	81 
    -- CP-element group 29: 	73 
    -- CP-element group 29: 	60 
    -- CP-element group 29: 	63 
    -- CP-element group 29: 	19 
    -- CP-element group 29: 	69 
    -- CP-element group 29: 	23 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (15) 
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_resized_1
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_computed_1
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_resize_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_resize_1/index_resize_req
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_resize_1/index_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_final_index_sum_regn_Sample/req
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_scale_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_scale_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_scale_1/scale_rename_req
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_scale_1/scale_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_resize_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_final_index_sum_regn_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_index_scaled_1
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_update_completed__ps
      -- 
    req_974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(29), ack => array_obj_ref_413_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	16 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_loopback_trigger
      -- 
    loadKernelChannel_CP_671_elements(30) <= loadKernelChannel_CP_671_elements(16);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_loopback_sample_req
      -- CP-element group 31: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_loopback_sample_req_ps
      -- 
    phi_stmt_363_loopback_sample_req_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_363_loopback_sample_req_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(31), ack => phi_stmt_363_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(31) is bound as output of CP function.
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_entry_trigger
      -- 
    loadKernelChannel_CP_671_elements(32) <= loadKernelChannel_CP_671_elements(17);
    -- CP-element group 33:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_entry_sample_req
      -- CP-element group 33: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_entry_sample_req_ps
      -- 
    phi_stmt_363_entry_sample_req_826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_363_entry_sample_req_826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(33), ack => phi_stmt_363_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_phi_mux_ack
      -- CP-element group 34: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_363_phi_mux_ack_ps
      -- 
    phi_stmt_363_phi_mux_ack_829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_363_ack_0, ack => loadKernelChannel_CP_671_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_Sample/req
      -- 
    req_842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(35), ack => nmycount_385_365_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_update_start__ps
      -- CP-element group 36: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_update_start_
      -- CP-element group 36: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_Update/req
      -- 
    req_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(36), ack => nmycount_385_365_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_sample_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_Sample/ack
      -- 
    ack_843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_385_365_buf_ack_0, ack => loadKernelChannel_CP_671_elements(37)); -- 
    -- CP-element group 38:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_update_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nmycount_365_Update/ack
      -- 
    ack_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_385_365_buf_ack_1, ack => loadKernelChannel_CP_671_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_sample_start__ps
      -- CP-element group 39: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_Sample/req
      -- 
    req_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(39), ack => start_add_366_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_Update/req
      -- CP-element group 40: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_update_start__ps
      -- CP-element group 40: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_update_start_
      -- CP-element group 40: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_Update/$entry
      -- 
    req_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(40), ack => start_add_366_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(40) is bound as output of CP function.
    -- CP-element group 41:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_sample_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_Sample/ack
      -- 
    ack_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_366_buf_ack_0, ack => loadKernelChannel_CP_671_elements(41)); -- 
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_update_completed__ps
      -- CP-element group 42: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_start_add_366_update_completed_
      -- 
    ack_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_366_buf_ack_1, ack => loadKernelChannel_CP_671_elements(42)); -- 
    -- CP-element group 43:  join  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	18 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	84 
    -- CP-element group 43: 	88 
    -- CP-element group 43: 	21 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	20 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_sample_start_
      -- 
    loadKernelChannel_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(80) & loadKernelChannel_CP_671_elements(84) & loadKernelChannel_CP_671_elements(88) & loadKernelChannel_CP_671_elements(21);
      gj_loadKernelChannel_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	18 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	87 
    -- CP-element group 44: 	46 
    -- CP-element group 44: 	61 
    -- CP-element group 44: 	64 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	22 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_update_start_
      -- 
    loadKernelChannel_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(87) & loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(61) & loadKernelChannel_CP_671_elements(64);
      gj_loadKernelChannel_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	21 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_671_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	85 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	63 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_update_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_671_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_loopback_trigger
      -- 
    loadKernelChannel_CP_671_elements(47) <= loadKernelChannel_CP_671_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_loopback_sample_req
      -- CP-element group 48: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_loopback_sample_req_ps
      -- 
    phi_stmt_367_loopback_sample_req_877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_367_loopback_sample_req_877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(48), ack => phi_stmt_367_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_entry_trigger
      -- 
    loadKernelChannel_CP_671_elements(49) <= loadKernelChannel_CP_671_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_entry_sample_req
      -- CP-element group 50: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_entry_sample_req_ps
      -- 
    phi_stmt_367_entry_sample_req_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_367_entry_sample_req_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(50), ack => phi_stmt_367_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_phi_mux_ack
      -- CP-element group 51: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/phi_stmt_367_phi_mux_ack_ps
      -- 
    phi_stmt_367_phi_mux_ack_883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_367_ack_0, ack => loadKernelChannel_CP_671_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_Sample/req
      -- 
    req_896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(52), ack => my_fetch_350_369_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_update_start_
      -- CP-element group 53: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_Update/req
      -- 
    req_901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(53), ack => my_fetch_350_369_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_Sample/ack
      -- 
    ack_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_350_369_buf_ack_0, ack => loadKernelChannel_CP_671_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_my_fetch_369_Update/ack
      -- 
    ack_902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_350_369_buf_ack_1, ack => loadKernelChannel_CP_671_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_sample_start_
      -- 
    req_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(56), ack => nfetch_val_435_370_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_update_start_
      -- CP-element group 57: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_Update/req
      -- CP-element group 57: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_update_start__ps
      -- 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(57), ack => nfetch_val_435_370_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_sample_completed__ps
      -- 
    ack_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_435_370_buf_ack_0, ack => loadKernelChannel_CP_671_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/R_nfetch_val_370_update_completed__ps
      -- 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_435_370_buf_ack_1, ack => loadKernelChannel_CP_671_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	46 
    -- CP-element group 60: 	29 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_Sample/$entry
      -- 
    req_929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(60), ack => WPIPE_kernel_pipe1_393_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(29) & loadKernelChannel_CP_671_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	44 
    -- CP-element group 61: 	25 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_update_start_
      -- CP-element group 61: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_Update/req
      -- 
    ack_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_393_inst_ack_0, ack => loadKernelChannel_CP_671_elements(61)); -- 
    req_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(61), ack => WPIPE_kernel_pipe1_393_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	90 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe1_393_Update/$exit
      -- 
    ack_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_393_inst_ack_1, ack => loadKernelChannel_CP_671_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	46 
    -- CP-element group 63: 	29 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_sample_start_
      -- 
    req_943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(63), ack => WPIPE_kernel_pipe2_397_inst_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(29) & loadKernelChannel_CP_671_elements(65);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	44 
    -- CP-element group 64: 	25 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_Update/req
      -- CP-element group 64: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_update_start_
      -- CP-element group 64: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_sample_completed_
      -- 
    ack_944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_397_inst_ack_0, ack => loadKernelChannel_CP_671_elements(64)); -- 
    req_948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(64), ack => WPIPE_kernel_pipe2_397_inst_req_1); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	90 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_Update/ack
      -- CP-element group 65: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/WPIPE_kernel_pipe2_397_update_completed_
      -- 
    ack_949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_397_inst_ack_1, ack => loadKernelChannel_CP_671_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	70 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	71 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	71 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_request/req
      -- CP-element group 66: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_request/$entry
      -- CP-element group 66: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_sample_start_
      -- 
    req_989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(66), ack => addr_of_414_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(70) & loadKernelChannel_CP_671_elements(71);
      gj_loadKernelChannel_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	18 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	72 
    -- CP-element group 67: 	79 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	72 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_update_start_
      -- CP-element group 67: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_complete/req
      -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(67), ack => addr_of_414_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(72) & loadKernelChannel_CP_671_elements(79);
      gj_loadKernelChannel_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	18 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: 	71 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_final_index_sum_regn_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_final_index_sum_regn_Update/req
      -- CP-element group 68: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_final_index_sum_regn_update_start
      -- 
    req_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(68), ack => array_obj_ref_413_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(70) & loadKernelChannel_CP_671_elements(71);
      gj_loadKernelChannel_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	29 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	90 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	25 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_final_index_sum_regn_Sample/ack
      -- CP-element group 69: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_final_index_sum_regn_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_final_index_sum_regn_sample_complete
      -- 
    ack_975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_413_index_offset_ack_0, ack => loadKernelChannel_CP_671_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	66 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (8) 
      -- CP-element group 70: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_final_index_sum_regn_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_offset_calculated
      -- CP-element group 70: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_final_index_sum_regn_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/array_obj_ref_413_root_address_calculated
      -- 
    ack_980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_413_index_offset_ack_1, ack => loadKernelChannel_CP_671_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	66 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	66 
    -- CP-element group 71: 	68 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_request/$exit
      -- CP-element group 71: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_request/ack
      -- 
    ack_990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_414_final_reg_ack_0, ack => loadKernelChannel_CP_671_elements(71)); -- 
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	67 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	77 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	67 
    -- CP-element group 72:  members (19) 
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_word_addrgen/root_register_ack
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_word_addrgen/$entry
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_word_addrgen/root_register_req
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_complete/$exit
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_complete/ack
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/addr_of_414_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_word_addrgen/$exit
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_base_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_base_plus_offset/$exit
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_base_plus_offset/$entry
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_base_addr_resize/base_resize_ack
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_base_addr_resize/base_resize_req
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_base_addr_resize/$exit
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_base_addr_resize/$entry
      -- CP-element group 72: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_base_address_resized
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_414_final_reg_ack_1, ack => loadKernelChannel_CP_671_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	29 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_Sample/req
      -- 
    req_1003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(73), ack => W_fn_404_delayed_7_0_416_inst_req_0); -- 
    loadKernelChannel_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(29) & loadKernelChannel_CP_671_elements(75);
      gj_loadKernelChannel_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: 	79 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_update_start_
      -- CP-element group 74: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_Update/req
      -- 
    req_1008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(74), ack => W_fn_404_delayed_7_0_416_inst_req_1); -- 
    loadKernelChannel_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(76) & loadKernelChannel_CP_671_elements(79);
      gj_loadKernelChannel_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	25 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_Sample/ack
      -- 
    ack_1004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_404_delayed_7_0_416_inst_ack_0, ack => loadKernelChannel_CP_671_elements(75)); -- 
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_Update/ack
      -- CP-element group 76: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_418_Update/$exit
      -- 
    ack_1009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_404_delayed_7_0_416_inst_ack_1, ack => loadKernelChannel_CP_671_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	72 
    -- CP-element group 77: 	76 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_sample_start_
      -- 
    rr_1042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(77), ack => ptr_deref_422_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(72) & loadKernelChannel_CP_671_elements(76) & loadKernelChannel_CP_671_elements(79);
      gj_loadKernelChannel_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	21 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_update_start_
      -- CP-element group 78: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/word_access_complete/$entry
      -- CP-element group 78: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/word_access_complete/word_0/$entry
      -- CP-element group 78: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/word_access_complete/word_0/cr
      -- 
    cr_1053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(78), ack => ptr_deref_422_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(80);
      gj_loadKernelChannel_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	74 
    -- CP-element group 79: 	77 
    -- CP-element group 79: 	67 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Sample/word_access_start/word_0/ra
      -- CP-element group 79: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Sample/word_access_start/$exit
      -- CP-element group 79: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Sample/word_access_start/word_0/$exit
      -- 
    ra_1043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_422_load_0_ack_0, ack => loadKernelChannel_CP_671_elements(79)); -- 
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	90 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	43 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/ptr_deref_422_Merge/merge_req
      -- CP-element group 80: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/ptr_deref_422_Merge/$exit
      -- CP-element group 80: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/ptr_deref_422_Merge/merge_ack
      -- CP-element group 80: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/word_access_complete/$exit
      -- CP-element group 80: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/word_access_complete/word_0/$exit
      -- CP-element group 80: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/word_access_complete/word_0/ca
      -- CP-element group 80: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/ptr_deref_422_Update/ptr_deref_422_Merge/$entry
      -- 
    ca_1054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_422_load_0_ack_1, ack => loadKernelChannel_CP_671_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	29 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_Sample/req
      -- CP-element group 81: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_sample_start_
      -- 
    req_1067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(81), ack => W_fn_410_delayed_13_0_424_inst_req_0); -- 
    loadKernelChannel_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(29) & loadKernelChannel_CP_671_elements(83);
      gj_loadKernelChannel_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	21 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_Update/req
      -- CP-element group 82: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_update_start_
      -- 
    req_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(82), ack => W_fn_410_delayed_13_0_424_inst_req_1); -- 
    loadKernelChannel_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(84);
      gj_loadKernelChannel_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	25 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_Sample/ack
      -- CP-element group 83: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_sample_completed_
      -- 
    ack_1068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_410_delayed_13_0_424_inst_ack_0, ack => loadKernelChannel_CP_671_elements(83)); -- 
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	90 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	43 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_Update/ack
      -- CP-element group 84: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_426_update_completed_
      -- 
    ack_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_410_delayed_13_0_424_inst_ack_1, ack => loadKernelChannel_CP_671_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	46 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_Sample/req
      -- 
    req_1081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(85), ack => W_fetch_val_412_delayed_13_0_427_inst_req_0); -- 
    loadKernelChannel_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(87);
      gj_loadKernelChannel_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	21 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_Update/req
      -- CP-element group 86: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_update_start_
      -- 
    req_1086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(86), ack => W_fetch_val_412_delayed_13_0_427_inst_req_1); -- 
    loadKernelChannel_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(88);
      gj_loadKernelChannel_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	44 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_sample_completed_
      -- 
    ack_1082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_412_delayed_13_0_427_inst_ack_0, ack => loadKernelChannel_CP_671_elements(87)); -- 
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	43 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/assign_stmt_429_update_completed_
      -- 
    ack_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_412_delayed_13_0_427_inst_ack_1, ack => loadKernelChannel_CP_671_elements(88)); -- 
    -- CP-element group 89:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	18 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	19 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_671_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_671_elements(18), ack => loadKernelChannel_CP_671_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	80 
    -- CP-element group 90: 	84 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	65 
    -- CP-element group 90: 	62 
    -- CP-element group 90: 	69 
    -- CP-element group 90: 	21 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	15 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_360/do_while_stmt_361/do_while_stmt_361_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(80) & loadKernelChannel_CP_671_elements(84) & loadKernelChannel_CP_671_elements(88) & loadKernelChannel_CP_671_elements(65) & loadKernelChannel_CP_671_elements(62) & loadKernelChannel_CP_671_elements(69) & loadKernelChannel_CP_671_elements(21);
      gj_loadKernelChannel_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	14 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_360/do_while_stmt_361/loop_exit/ack
      -- CP-element group 91: 	 branch_block_stmt_360/do_while_stmt_361/loop_exit/$exit
      -- 
    ack_1092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_361_branch_ack_0, ack => loadKernelChannel_CP_671_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	14 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_360/do_while_stmt_361/loop_taken/$exit
      -- CP-element group 92: 	 branch_block_stmt_360/do_while_stmt_361/loop_taken/ack
      -- 
    ack_1096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_361_branch_ack_1, ack => loadKernelChannel_CP_671_elements(92)); -- 
    -- CP-element group 93:  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	12 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	10 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_360/do_while_stmt_361/$exit
      -- 
    loadKernelChannel_CP_671_elements(93) <= loadKernelChannel_CP_671_elements(12);
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	10 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 assign_stmt_451/CONCAT_u1_u32_450_Sample/ra
      -- CP-element group 94: 	 assign_stmt_451/CONCAT_u1_u32_450_Sample/$exit
      -- CP-element group 94: 	 assign_stmt_451/CONCAT_u1_u32_450_sample_completed_
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u32_450_inst_ack_0, ack => loadKernelChannel_CP_671_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	10 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 assign_stmt_451/WPIPE_size_pipe_443_Sample/req
      -- CP-element group 95: 	 assign_stmt_451/CONCAT_u1_u32_450_Update/ca
      -- CP-element group 95: 	 assign_stmt_451/WPIPE_size_pipe_443_sample_start_
      -- CP-element group 95: 	 assign_stmt_451/CONCAT_u1_u32_450_update_completed_
      -- CP-element group 95: 	 assign_stmt_451/WPIPE_size_pipe_443_Sample/$entry
      -- CP-element group 95: 	 assign_stmt_451/CONCAT_u1_u32_450_Update/$exit
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u32_450_inst_ack_1, ack => loadKernelChannel_CP_671_elements(95)); -- 
    req_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(95), ack => WPIPE_size_pipe_443_inst_req_0); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (6) 
      -- CP-element group 96: 	 assign_stmt_451/WPIPE_size_pipe_443_Sample/ack
      -- CP-element group 96: 	 assign_stmt_451/WPIPE_size_pipe_443_Update/$entry
      -- CP-element group 96: 	 assign_stmt_451/WPIPE_size_pipe_443_Update/req
      -- CP-element group 96: 	 assign_stmt_451/WPIPE_size_pipe_443_sample_completed_
      -- CP-element group 96: 	 assign_stmt_451/WPIPE_size_pipe_443_update_start_
      -- CP-element group 96: 	 assign_stmt_451/WPIPE_size_pipe_443_Sample/$exit
      -- 
    ack_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_443_inst_ack_0, ack => loadKernelChannel_CP_671_elements(96)); -- 
    req_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(96), ack => WPIPE_size_pipe_443_inst_req_1); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 assign_stmt_451/$exit
      -- CP-element group 97: 	 assign_stmt_451/WPIPE_size_pipe_443_Update/$exit
      -- CP-element group 97: 	 assign_stmt_451/WPIPE_size_pipe_443_Update/ack
      -- CP-element group 97: 	 assign_stmt_451/WPIPE_size_pipe_443_update_completed_
      -- CP-element group 97: 	 $exit
      -- 
    ack_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_443_inst_ack_1, ack => loadKernelChannel_CP_671_elements(97)); -- 
    loadKernelChannel_do_while_stmt_361_terminator_1097: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_361_terminator_1097", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_671_elements(15),loop_continue => loadKernelChannel_CP_671_elements(92),loop_terminate => loadKernelChannel_CP_671_elements(91),loop_back => loadKernelChannel_CP_671_elements(13),loop_exit => loadKernelChannel_CP_671_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_363_phi_seq_867_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_671_elements(30);
      loadKernelChannel_CP_671_elements(35)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_671_elements(37);
      loadKernelChannel_CP_671_elements(36)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_671_elements(38);
      loadKernelChannel_CP_671_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_671_elements(32);
      loadKernelChannel_CP_671_elements(39)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_671_elements(41);
      loadKernelChannel_CP_671_elements(40)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_671_elements(42);
      loadKernelChannel_CP_671_elements(33) <= phi_mux_reqs(1);
      phi_stmt_363_phi_seq_867 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_363_phi_seq_867") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_671_elements(26), 
          phi_sample_ack => loadKernelChannel_CP_671_elements(27), 
          phi_update_req => loadKernelChannel_CP_671_elements(28), 
          phi_update_ack => loadKernelChannel_CP_671_elements(29), 
          phi_mux_ack => loadKernelChannel_CP_671_elements(34), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_367_phi_seq_921_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_671_elements(49);
      loadKernelChannel_CP_671_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_671_elements(54);
      loadKernelChannel_CP_671_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_671_elements(55);
      loadKernelChannel_CP_671_elements(50) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_671_elements(47);
      loadKernelChannel_CP_671_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_671_elements(58);
      loadKernelChannel_CP_671_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_671_elements(59);
      loadKernelChannel_CP_671_elements(48) <= phi_mux_reqs(1);
      phi_stmt_367_phi_seq_921 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_367_phi_seq_921") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_671_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_671_elements(45), 
          phi_update_req => loadKernelChannel_CP_671_elements(22), 
          phi_update_ack => loadKernelChannel_CP_671_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_671_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_809_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_671_elements(16);
        preds(1)  <= loadKernelChannel_CP_671_elements(17);
        entry_tmerge_809 : transition_merge -- 
          generic map(name => " entry_tmerge_809")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_671_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_376_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_403_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u1_u32_450_wire : std_logic_vector(31 downto 0);
    signal LSHR_u64_u64_389_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_412_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_412_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_412_wire : std_logic_vector(63 downto 0);
    signal R_sh_start_343_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_343_scaled : std_logic_vector(13 downto 0);
    signal SUB_u64_u64_377_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_440_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_448_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_441_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_344_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_344_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_344_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_344_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_344_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_344_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_413_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_413_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_413_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_413_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_413_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_413_root_address : std_logic_vector(13 downto 0);
    signal fetch_addr_346 : std_logic_vector(31 downto 0);
    signal fetch_addr_415 : std_logic_vector(31 downto 0);
    signal fetch_val_367 : std_logic_vector(63 downto 0);
    signal fetch_val_412_delayed_13_0_429 : std_logic_vector(63 downto 0);
    signal first_fill_355 : std_logic_vector(0 downto 0);
    signal fn_404_delayed_7_0_418 : std_logic_vector(0 downto 0);
    signal fn_406 : std_logic_vector(0 downto 0);
    signal fn_410_delayed_13_0_426 : std_logic_vector(0 downto 0);
    signal fv_423 : std_logic_vector(63 downto 0);
    signal konst_333_wire_constant : std_logic_vector(63 downto 0);
    signal konst_353_wire_constant : std_logic_vector(63 downto 0);
    signal konst_373_wire_constant : std_logic_vector(63 downto 0);
    signal konst_375_wire_constant : std_logic_vector(63 downto 0);
    signal konst_378_wire_constant : std_logic_vector(63 downto 0);
    signal konst_383_wire_constant : std_logic_vector(63 downto 0);
    signal konst_402_wire_constant : std_logic_vector(63 downto 0);
    signal konst_404_wire_constant : std_logic_vector(63 downto 0);
    signal konst_411_wire_constant : std_logic_vector(63 downto 0);
    signal konst_439_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_350 : std_logic_vector(63 downto 0);
    signal my_fetch_350_369_buffered : std_logic_vector(63 downto 0);
    signal my_num1_380 : std_logic_vector(63 downto 0);
    signal mycount_363 : std_logic_vector(63 downto 0);
    signal nfetch_val_435 : std_logic_vector(63 downto 0);
    signal nfetch_val_435_370_buffered : std_logic_vector(63 downto 0);
    signal nmycount_385 : std_logic_vector(63 downto 0);
    signal nmycount_385_365_buffered : std_logic_vector(63 downto 0);
    signal pingpong_339 : std_logic_vector(0 downto 0);
    signal ptr_deref_349_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_349_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_349_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_349_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_349_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_422_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_422_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_422_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_422_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_422_word_offset_0 : std_logic_vector(13 downto 0);
    signal sh_start_335 : std_logic_vector(63 downto 0);
    signal start_add_366_buffered : std_logic_vector(63 downto 0);
    signal start_next_359 : std_logic_vector(0 downto 0);
    signal type_cast_449_wire : std_logic_vector(30 downto 0);
    signal var_val_391 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_344_constant_part_of_offset <= "00000000000000";
    array_obj_ref_344_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_344_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_344_resized_base_address <= "00000000000000";
    array_obj_ref_413_constant_part_of_offset <= "00000000000000";
    array_obj_ref_413_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_413_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_413_resized_base_address <= "00000000000000";
    konst_333_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_353_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_373_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_375_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_378_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_383_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_402_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_404_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_411_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_439_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_349_word_offset_0 <= "00000000000000";
    ptr_deref_422_word_offset_0 <= "00000000000000";
    phi_stmt_363: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_385_365_buffered & start_add_366_buffered;
      req <= phi_stmt_363_req_0 & phi_stmt_363_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_363",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_363_ack_0,
          idata => idata,
          odata => mycount_363,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_363
    phi_stmt_367: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch_350_369_buffered & nfetch_val_435_370_buffered;
      req <= phi_stmt_367_req_0 & phi_stmt_367_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_367",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_367_ack_0,
          idata => idata,
          odata => fetch_val_367,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_367
    -- flow-through select operator MUX_434_inst
    nfetch_val_435 <= fv_423 when (fn_410_delayed_13_0_426(0) /=  '0') else fetch_val_412_delayed_13_0_429;
    W_fetch_val_412_delayed_13_0_427_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_412_delayed_13_0_427_inst_req_0;
      W_fetch_val_412_delayed_13_0_427_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_412_delayed_13_0_427_inst_req_1;
      W_fetch_val_412_delayed_13_0_427_inst_ack_1<= rack(0);
      W_fetch_val_412_delayed_13_0_427_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_412_delayed_13_0_427_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_412_delayed_13_0_429,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_404_delayed_7_0_416_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_404_delayed_7_0_416_inst_req_0;
      W_fn_404_delayed_7_0_416_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_404_delayed_7_0_416_inst_req_1;
      W_fn_404_delayed_7_0_416_inst_ack_1<= rack(0);
      W_fn_404_delayed_7_0_416_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_404_delayed_7_0_416_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_404_delayed_7_0_418,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_410_delayed_13_0_424_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_410_delayed_13_0_424_inst_req_0;
      W_fn_410_delayed_13_0_424_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_410_delayed_13_0_424_inst_req_1;
      W_fn_410_delayed_13_0_424_inst_ack_1<= rack(0);
      W_fn_410_delayed_13_0_424_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_410_delayed_13_0_424_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_410_delayed_13_0_426,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_345_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_345_final_reg_req_0;
      addr_of_345_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_345_final_reg_req_1;
      addr_of_345_final_reg_ack_1<= rack(0);
      addr_of_345_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_345_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_344_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_414_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_414_final_reg_req_0;
      addr_of_414_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_414_final_reg_req_1;
      addr_of_414_final_reg_ack_1<= rack(0);
      addr_of_414_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_414_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_413_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_415,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_350_369_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_350_369_buf_req_0;
      my_fetch_350_369_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_350_369_buf_req_1;
      my_fetch_350_369_buf_ack_1<= rack(0);
      my_fetch_350_369_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_350_369_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_350,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_350_369_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_435_370_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_435_370_buf_req_0;
      nfetch_val_435_370_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_435_370_buf_req_1;
      nfetch_val_435_370_buf_ack_1<= rack(0);
      nfetch_val_435_370_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_435_370_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_435,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_435_370_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_385_365_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_385_365_buf_req_0;
      nmycount_385_365_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_385_365_buf_req_1;
      nmycount_385_365_buf_ack_1<= rack(0);
      nmycount_385_365_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_385_365_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_385_365_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_366_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_366_buf_req_0;
      start_add_366_buf_ack_0<= wack(0);
      rreq(0) <= start_add_366_buf_req_1;
      start_add_366_buf_ack_1<= rack(0);
      start_add_366_buf : InterlockBuffer generic map ( -- 
        name => "start_add_366_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_366_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_338_inst
    process(pp_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := pp_buffer(0 downto 0);
      pingpong_339 <= tmp_var; -- 
    end process;
    -- interlock type_cast_390_inst
    process(LSHR_u64_u64_389_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_389_wire(15 downto 0);
      var_val_391 <= tmp_var; -- 
    end process;
    -- interlock type_cast_449_inst
    process(SUB_u64_u64_448_wire) -- 
      variable tmp_var : std_logic_vector(30 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 30 downto 0) := SUB_u64_u64_448_wire(30 downto 0);
      type_cast_449_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_344_index_1_rename
    process(R_sh_start_343_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_343_resized;
      ov(13 downto 0) := iv;
      R_sh_start_343_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_344_index_1_resize
    process(sh_start_335) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_335;
      ov := iv(13 downto 0);
      R_sh_start_343_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_344_root_address_inst
    process(array_obj_ref_344_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_344_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_344_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_413_index_1_rename
    process(LSHR_u64_u64_412_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_412_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_412_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_413_index_1_resize
    process(LSHR_u64_u64_412_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_412_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_412_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_413_root_address_inst
    process(array_obj_ref_413_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_413_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_413_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_addr_0
    process(ptr_deref_349_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_349_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_349_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_base_resize
    process(fetch_addr_346) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_346;
      ov := iv(13 downto 0);
      ptr_deref_349_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_gather_scatter
    process(ptr_deref_349_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_349_data_0;
      ov(63 downto 0) := iv;
      my_fetch_350 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_root_address_inst
    process(ptr_deref_349_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_349_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_349_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_422_addr_0
    process(ptr_deref_422_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_422_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_422_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_422_base_resize
    process(fetch_addr_415) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_415;
      ov := iv(13 downto 0);
      ptr_deref_422_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_422_gather_scatter
    process(ptr_deref_422_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_422_data_0;
      ov(63 downto 0) := iv;
      fv_423 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_422_root_address_inst
    process(ptr_deref_422_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_422_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_422_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_361_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_441_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_361_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_361_branch_req_0,
          ack0 => do_while_stmt_361_branch_ack_0,
          ack1 => do_while_stmt_361_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_384_inst
    process(mycount_363) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_363, konst_383_wire_constant, tmp_var);
      nmycount_385 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_376_inst
    process(mycount_363) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_363, konst_375_wire_constant, tmp_var);
      AND_u64_u64_376_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_403_inst
    process(nmycount_385) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_385, konst_402_wire_constant, tmp_var);
      AND_u64_u64_403_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : CONCAT_u1_u32_450_inst 
    ApConcat_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pingpong_339 & type_cast_449_wire;
      CONCAT_u1_u32_450_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u1_u32_450_inst_req_0;
      CONCAT_u1_u32_450_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u1_u32_450_inst_req_1;
      CONCAT_u1_u32_450_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_3_gI: SplitGuardInterface generic map(name => "ApConcat_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 31, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- binary operator EQ_u64_u1_354_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_353_wire_constant, tmp_var);
      first_fill_355 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_405_inst
    process(AND_u64_u64_403_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_403_wire, konst_404_wire_constant, tmp_var);
      fn_406 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_334_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_333_wire_constant, tmp_var);
      sh_start_335 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_389_inst
    process(fetch_val_367, my_num1_380) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_367, my_num1_380, tmp_var);
      LSHR_u64_u64_389_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_412_inst
    process(nmycount_385) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_385, konst_411_wire_constant, tmp_var);
      LSHR_u64_u64_412_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_379_inst
    process(SUB_u64_u64_377_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_377_wire, konst_378_wire_constant, tmp_var);
      my_num1_380 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_377_inst
    process(konst_373_wire_constant, AND_u64_u64_376_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_373_wire_constant, AND_u64_u64_376_wire, tmp_var);
      SUB_u64_u64_377_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_440_inst
    process(end_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, konst_439_wire_constant, tmp_var);
      SUB_u64_u64_440_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_448_inst
    process(end_add_buffer, start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, start_add_buffer, tmp_var);
      SUB_u64_u64_448_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_441_inst
    process(mycount_363, SUB_u64_u64_440_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_363, SUB_u64_u64_440_wire, tmp_var);
      ULT_u64_u1_441_wire <= tmp_var; --
    end process;
    -- shared split operator group (14) : array_obj_ref_344_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_343_scaled;
      array_obj_ref_344_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_344_index_offset_req_0;
      array_obj_ref_344_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_344_index_offset_req_1;
      array_obj_ref_344_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : array_obj_ref_413_index_offset 
    ApIntAdd_group_15: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_412_scaled;
      array_obj_ref_413_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_413_index_offset_req_0;
      array_obj_ref_413_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_413_index_offset_req_1;
      array_obj_ref_413_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_15_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared load operator group (0) : ptr_deref_349_load_0 ptr_deref_422_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_349_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_422_load_0_req_0;
      ptr_deref_349_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_422_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_349_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_422_load_0_req_1;
      ptr_deref_349_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_422_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_404_delayed_7_0_418(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_349_word_address_0 & ptr_deref_422_word_address_0;
      ptr_deref_349_data_0 <= data_out(127 downto 64);
      ptr_deref_422_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_358_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_358_inst_req_0;
      RPIPE_input_done_pipe_358_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_358_inst_req_1;
      RPIPE_input_done_pipe_358_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_355(0);
      start_next_359 <= data_out(0 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_393_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_393_inst_req_0;
      WPIPE_kernel_pipe1_393_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_393_inst_req_1;
      WPIPE_kernel_pipe1_393_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  not pingpong_339(0);
      data_in <= var_val_391;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe2_397_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe2_397_inst_req_0;
      WPIPE_kernel_pipe2_397_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe2_397_inst_req_1;
      WPIPE_kernel_pipe2_397_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= pingpong_339(0);
      data_in <= var_val_391;
      kernel_pipe2_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe2_pipe_write_req(0),
          oack => kernel_pipe2_pipe_write_ack(0),
          odata => kernel_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_size_pipe_443_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_443_inst_req_0;
      WPIPE_size_pipe_443_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_443_inst_req_1;
      WPIPE_size_pipe_443_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u1_u32_450_wire;
      size_pipe_write_2_gI: SplitGuardInterface generic map(name => "size_pipe_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_637_start: Boolean;
  signal timer_CP_637_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_319_inst_req_0 : boolean;
  signal WPIPE_timer_req_319_inst_ack_0 : boolean;
  signal WPIPE_timer_req_319_inst_req_1 : boolean;
  signal WPIPE_timer_req_319_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_324_inst_req_0 : boolean;
  signal RPIPE_timer_resp_324_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_324_inst_req_1 : boolean;
  signal RPIPE_timer_resp_324_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_637_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_637: Block -- control-path 
    signal timer_CP_637_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_637_elements(0) <= timer_CP_637_start;
    timer_CP_637_symbol <= timer_CP_637_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_322_to_assign_stmt_325/$entry
      -- CP-element group 0: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_sample_start_
      -- CP-element group 0: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_Sample/req
      -- CP-element group 0: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_sample_start_
      -- CP-element group 0: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_Sample/rr
      -- 
    req_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => WPIPE_timer_req_319_inst_req_0); -- 
    rr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => RPIPE_timer_resp_324_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_sample_completed_
      -- CP-element group 1: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_update_start_
      -- CP-element group 1: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_Sample/ack
      -- CP-element group 1: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_Update/$entry
      -- CP-element group 1: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_Update/req
      -- 
    ack_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_319_inst_ack_0, ack => timer_CP_637_elements(1)); -- 
    req_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(1), ack => WPIPE_timer_req_319_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_update_completed_
      -- CP-element group 2: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_Update/$exit
      -- CP-element group 2: 	 assign_stmt_322_to_assign_stmt_325/WPIPE_timer_req_319_Update/ack
      -- 
    ack_656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_319_inst_ack_1, ack => timer_CP_637_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_sample_completed_
      -- CP-element group 3: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_update_start_
      -- CP-element group 3: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_Sample/ra
      -- CP-element group 3: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_Update/$entry
      -- CP-element group 3: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_Update/cr
      -- 
    ra_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_324_inst_ack_0, ack => timer_CP_637_elements(3)); -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(3), ack => RPIPE_timer_resp_324_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_update_completed_
      -- CP-element group 4: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_Update/$exit
      -- CP-element group 4: 	 assign_stmt_322_to_assign_stmt_325/RPIPE_timer_resp_324_Update/ca
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_324_inst_ack_1, ack => timer_CP_637_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_322_to_assign_stmt_325/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_637_elements(2) & timer_CP_637_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_637_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_321_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_321_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_324_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_324_inst_req_0;
      RPIPE_timer_resp_324_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_324_inst_req_1;
      RPIPE_timer_resp_324_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_319_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_319_inst_req_0;
      WPIPE_timer_req_319_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_319_inst_req_1;
      WPIPE_timer_req_319_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_321_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_4687_start: Boolean;
  signal timerDaemon_CP_4687_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_2073_branch_ack_0 : boolean;
  signal RPIPE_timer_req_2082_inst_req_0 : boolean;
  signal RPIPE_timer_req_2082_inst_ack_0 : boolean;
  signal RPIPE_timer_req_2082_inst_req_1 : boolean;
  signal RPIPE_timer_req_2082_inst_ack_1 : boolean;
  signal do_while_stmt_2073_branch_ack_1 : boolean;
  signal WPIPE_timer_resp_2090_inst_req_0 : boolean;
  signal WPIPE_timer_resp_2090_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_2090_inst_req_1 : boolean;
  signal phi_stmt_2075_ack_0 : boolean;
  signal nCOUNTER_2088_2079_buf_ack_1 : boolean;
  signal nCOUNTER_2088_2079_buf_req_1 : boolean;
  signal phi_stmt_2075_req_0 : boolean;
  signal phi_stmt_2075_req_1 : boolean;
  signal nCOUNTER_2088_2079_buf_ack_0 : boolean;
  signal nCOUNTER_2088_2079_buf_req_0 : boolean;
  signal do_while_stmt_2073_branch_req_0 : boolean;
  signal WPIPE_timer_resp_2090_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_4687_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4687_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_4687_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4687_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_4687: Block -- control-path 
    signal timerDaemon_CP_4687_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_4687_elements(0) <= timerDaemon_CP_4687_start;
    timerDaemon_CP_4687_symbol <= timerDaemon_CP_4687_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_2072/do_while_stmt_2073__entry__
      -- CP-element group 0: 	 branch_block_stmt_2072/$entry
      -- CP-element group 0: 	 branch_block_stmt_2072/branch_block_stmt_2072__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_2072/do_while_stmt_2073__exit__
      -- CP-element group 1: 	 branch_block_stmt_2072/branch_block_stmt_2072__exit__
      -- CP-element group 1: 	 branch_block_stmt_2072/$exit
      -- CP-element group 1: 	 $exit
      -- 
    timerDaemon_CP_4687_elements(1) <= timerDaemon_CP_4687_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073__entry__
      -- CP-element group 2: 	 branch_block_stmt_2072/do_while_stmt_2073/$entry
      -- 
    timerDaemon_CP_4687_elements(2) <= timerDaemon_CP_4687_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073__exit__
      -- 
    -- Element group timerDaemon_CP_4687_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2072/do_while_stmt_2073/loop_back
      -- 
    -- Element group timerDaemon_CP_4687_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2072/do_while_stmt_2073/condition_done
      -- CP-element group 5: 	 branch_block_stmt_2072/do_while_stmt_2073/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_2072/do_while_stmt_2073/loop_exit/$entry
      -- 
    timerDaemon_CP_4687_elements(5) <= timerDaemon_CP_4687_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2072/do_while_stmt_2073/loop_body_done
      -- 
    timerDaemon_CP_4687_elements(6) <= timerDaemon_CP_4687_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_4687_elements(7) <= timerDaemon_CP_4687_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_4687_elements(8) <= timerDaemon_CP_4687_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	32 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2080_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/$entry
      -- 
    -- Element group timerDaemon_CP_4687_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	40 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/condition_evaluated
      -- 
    condition_evaluated_4711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4687_elements(10), ack => do_while_stmt_2073_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(14) & timerDaemon_CP_4687_elements(40);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(9) & timerDaemon_CP_4687_elements(15) & timerDaemon_CP_4687_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2080_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/aggregated_phi_sample_ack
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(17) & timerDaemon_CP_4687_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(16) & timerDaemon_CP_4687_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(18) & timerDaemon_CP_4687_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(9) & timerDaemon_CP_4687_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(9) & timerDaemon_CP_4687_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_4687_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_4687_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_loopback_trigger
      -- 
    timerDaemon_CP_4687_elements(19) <= timerDaemon_CP_4687_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_loopback_sample_req
      -- 
    phi_stmt_2075_loopback_sample_req_4726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2075_loopback_sample_req_4726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4687_elements(20), ack => phi_stmt_2075_req_1); -- 
    -- Element group timerDaemon_CP_4687_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_entry_trigger
      -- 
    timerDaemon_CP_4687_elements(21) <= timerDaemon_CP_4687_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_entry_sample_req
      -- 
    phi_stmt_2075_entry_sample_req_4729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2075_entry_sample_req_4729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4687_elements(22), ack => phi_stmt_2075_req_0); -- 
    -- Element group timerDaemon_CP_4687_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2075_phi_mux_ack
      -- 
    phi_stmt_2075_phi_mux_ack_4732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2075_ack_0, ack => timerDaemon_CP_4687_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/type_cast_2078_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/type_cast_2078_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/type_cast_2078_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/type_cast_2078_sample_completed_
      -- 
    -- Element group timerDaemon_CP_4687_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/type_cast_2078_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/type_cast_2078_update_start_
      -- 
    -- Element group timerDaemon_CP_4687_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/type_cast_2078_update_completed__ps
      -- 
    timerDaemon_CP_4687_elements(26) <= timerDaemon_CP_4687_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/type_cast_2078_update_completed_
      -- 
    -- Element group timerDaemon_CP_4687_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_4687_elements(25), ack => timerDaemon_CP_4687_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_Sample/$entry
      -- 
    req_4753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4687_elements(28), ack => nCOUNTER_2088_2079_buf_req_0); -- 
    -- Element group timerDaemon_CP_4687_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_update_start_
      -- CP-element group 29: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_Update/req
      -- CP-element group 29: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_update_start__ps
      -- 
    req_4758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4687_elements(29), ack => nCOUNTER_2088_2079_buf_req_1); -- 
    -- Element group timerDaemon_CP_4687_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_Sample/$exit
      -- 
    ack_4754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_2088_2079_buf_ack_0, ack => timerDaemon_CP_4687_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/R_nCOUNTER_2079_update_completed_
      -- 
    ack_4759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_2088_2079_buf_ack_1, ack => timerDaemon_CP_4687_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2080_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(9) & timerDaemon_CP_4687_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_Sample/rr
      -- 
    rr_4772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4687_elements(33), ack => RPIPE_timer_req_2082_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(11) & timerDaemon_CP_4687_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_Update/cr
      -- 
    cr_4777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4687_elements(34), ack => RPIPE_timer_req_2082_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(13) & timerDaemon_CP_4687_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_Sample/$exit
      -- 
    ra_4773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_2082_inst_ack_0, ack => timerDaemon_CP_4687_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/phi_stmt_2080_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/RPIPE_timer_req_2082_Update/ca
      -- 
    ca_4778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_2082_inst_ack_1, ack => timerDaemon_CP_4687_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_Sample/req
      -- 
    req_4786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4687_elements(37), ack => WPIPE_timer_resp_2090_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(18) & timerDaemon_CP_4687_elements(36) & timerDaemon_CP_4687_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_update_start_
      -- CP-element group 38: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_Update/req
      -- 
    ack_4787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_2090_inst_ack_0, ack => timerDaemon_CP_4687_elements(38)); -- 
    req_4791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4687_elements(38), ack => WPIPE_timer_resp_2090_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/WPIPE_timer_resp_2090_Update/ack
      -- 
    ack_4792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_2090_inst_ack_1, ack => timerDaemon_CP_4687_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_4687_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_4687_elements(9), ack => timerDaemon_CP_4687_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2072/do_while_stmt_2073/do_while_stmt_2073_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4687_elements(12) & timerDaemon_CP_4687_elements(39);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4687_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_2072/do_while_stmt_2073/loop_exit/ack
      -- CP-element group 42: 	 branch_block_stmt_2072/do_while_stmt_2073/loop_exit/$exit
      -- 
    ack_4797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2073_branch_ack_0, ack => timerDaemon_CP_4687_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_2072/do_while_stmt_2073/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_2072/do_while_stmt_2073/loop_taken/ack
      -- 
    ack_4801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2073_branch_ack_1, ack => timerDaemon_CP_4687_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_2072/do_while_stmt_2073/$exit
      -- 
    timerDaemon_CP_4687_elements(44) <= timerDaemon_CP_4687_elements(3);
    timerDaemon_do_while_stmt_2073_terminator_4802: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_2073_terminator_4802", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_4687_elements(6),loop_continue => timerDaemon_CP_4687_elements(43),loop_terminate => timerDaemon_CP_4687_elements(42),loop_back => timerDaemon_CP_4687_elements(4),loop_exit => timerDaemon_CP_4687_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2075_phi_seq_4760_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_4687_elements(21);
      timerDaemon_CP_4687_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_4687_elements(24);
      timerDaemon_CP_4687_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_4687_elements(26);
      timerDaemon_CP_4687_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_4687_elements(19);
      timerDaemon_CP_4687_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_4687_elements(30);
      timerDaemon_CP_4687_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_4687_elements(31);
      timerDaemon_CP_4687_elements(20) <= phi_mux_reqs(1);
      phi_stmt_2075_phi_seq_4760 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_2075_phi_seq_4760") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_4687_elements(11), 
          phi_sample_ack => timerDaemon_CP_4687_elements(17), 
          phi_update_req => timerDaemon_CP_4687_elements(13), 
          phi_update_ack => timerDaemon_CP_4687_elements(18), 
          phi_mux_ack => timerDaemon_CP_4687_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4712_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_4687_elements(7);
        preds(1)  <= timerDaemon_CP_4687_elements(8);
        entry_tmerge_4712 : transition_merge -- 
          generic map(name => " entry_tmerge_4712")
          port map (preds => preds, symbol_out => timerDaemon_CP_4687_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_2075 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_2082_wire : std_logic_vector(0 downto 0);
    signal konst_2086_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2094_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_2088 : std_logic_vector(63 downto 0);
    signal nCOUNTER_2088_2079_buffered : std_logic_vector(63 downto 0);
    signal req_2080 : std_logic_vector(0 downto 0);
    signal type_cast_2078_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_2086_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_2094_wire_constant <= "1";
    type_cast_2078_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_2075: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2078_wire_constant & nCOUNTER_2088_2079_buffered;
      req <= phi_stmt_2075_req_0 & phi_stmt_2075_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2075",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2075_ack_0,
          idata => idata,
          odata => COUNTER_2075,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2075
    nCOUNTER_2088_2079_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_2088_2079_buf_req_0;
      nCOUNTER_2088_2079_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_2088_2079_buf_req_1;
      nCOUNTER_2088_2079_buf_ack_1<= rack(0);
      nCOUNTER_2088_2079_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_2088_2079_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_2088,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_2088_2079_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_2080
    process(RPIPE_timer_req_2082_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_2082_wire(0 downto 0);
      req_2080 <= tmp_var; -- 
    end process;
    do_while_stmt_2073_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2094_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2073_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2073_branch_req_0,
          ack0 => do_while_stmt_2073_branch_ack_0,
          ack1 => do_while_stmt_2073_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_2087_inst
    process(COUNTER_2075) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_2075, konst_2086_wire_constant, tmp_var);
      nCOUNTER_2088 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_2082_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_2082_inst_req_0;
      RPIPE_timer_req_2082_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_2082_inst_req_1;
      RPIPE_timer_req_2082_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_2082_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_2090_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_2090_inst_req_0;
      WPIPE_timer_resp_2090_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_2090_inst_req_1;
      WPIPE_timer_resp_2090_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_2080(0);
      data_in <= COUNTER_2075;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_num_cont :  std_logic_vector(15 downto 0);
  signal access_T_row1 :  std_logic_vector(15 downto 0);
  signal access_T_col1 :  std_logic_vector(15 downto 0);
  signal access_T_rk1 :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(95 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(95 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(95 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(135 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      pp : in  std_logic_vector(7 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_end_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_pp :  std_logic_vector(7 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(135 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(135 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(31 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(1 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe2
  signal kernel_pipe2_pipe_write_data: std_logic_vector(31 downto 0);
  signal kernel_pipe2_pipe_write_req: std_logic_vector(1 downto 0);
  signal kernel_pipe2_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe kernel_pipe2
  signal kernel_pipe2_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_num_cont <= access_T_in_args(95 downto 80);
  access_T_row1 <= access_T_in_args(79 downto 64);
  access_T_col1 <= access_T_in_args(63 downto 48);
  access_T_rk1 <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 96,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      num_cont => access_T_num_cont,
      row1 => access_T_row1,
      col1 => access_T_col1,
      rk1 => access_T_rk1,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(95 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(135 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      kernel_pipe2_pipe_read_req => kernel_pipe2_pipe_read_req(0 downto 0),
      kernel_pipe2_pipe_read_ack => kernel_pipe2_pipe_read_ack(0 downto 0),
      kernel_pipe2_pipe_read_data => kernel_pipe2_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(31 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(0 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      kernel_pipe2_pipe_write_req => kernel_pipe2_pipe_write_req(0 downto 0),
      kernel_pipe2_pipe_write_ack => kernel_pipe2_pipe_write_ack(0 downto 0),
      kernel_pipe2_pipe_write_data => kernel_pipe2_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(135 downto 72);
  loadKernelChannel_end_add <= loadKernelChannel_in_args(71 downto 8);
  loadKernelChannel_pp <= loadKernelChannel_in_args(7 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 136,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      end_add => loadKernelChannel_end_add,
      pp => loadKernelChannel_pp,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(0 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(1 downto 1),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(1 downto 1),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(31 downto 16),
      kernel_pipe2_pipe_write_req => kernel_pipe2_pipe_write_req(1 downto 1),
      kernel_pipe2_pipe_write_ack => kernel_pipe2_pipe_write_ack(1 downto 1),
      kernel_pipe2_pipe_write_data => kernel_pipe2_pipe_write_data(31 downto 16),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(31 downto 0),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe2",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => kernel_pipe2_pipe_read_req,
      read_ack => kernel_pipe2_pipe_read_ack,
      read_data => kernel_pipe2_pipe_read_data,
      write_req => kernel_pipe2_pipe_write_req,
      write_ack => kernel_pipe2_pipe_write_ack,
      write_data => kernel_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
