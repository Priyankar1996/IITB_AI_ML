-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendOutput_CP_26_start: Boolean;
  signal sendOutput_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_51_branch_req_0 : boolean;
  signal ptr_deref_81_load_0_req_1 : boolean;
  signal ptr_deref_81_load_0_ack_1 : boolean;
  signal if_stmt_51_branch_ack_1 : boolean;
  signal if_stmt_51_branch_ack_0 : boolean;
  signal type_cast_60_inst_req_0 : boolean;
  signal type_cast_60_inst_ack_0 : boolean;
  signal type_cast_60_inst_req_1 : boolean;
  signal type_cast_60_inst_ack_1 : boolean;
  signal array_obj_ref_76_index_offset_req_0 : boolean;
  signal array_obj_ref_76_index_offset_ack_0 : boolean;
  signal array_obj_ref_76_index_offset_req_1 : boolean;
  signal array_obj_ref_76_index_offset_ack_1 : boolean;
  signal addr_of_77_final_reg_req_0 : boolean;
  signal addr_of_77_final_reg_ack_0 : boolean;
  signal addr_of_77_final_reg_req_1 : boolean;
  signal addr_of_77_final_reg_ack_1 : boolean;
  signal ptr_deref_81_load_0_req_0 : boolean;
  signal ptr_deref_81_load_0_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_172_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_172_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_172_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_172_inst_ack_1 : boolean;
  signal type_cast_85_inst_req_0 : boolean;
  signal type_cast_85_inst_ack_0 : boolean;
  signal type_cast_85_inst_req_1 : boolean;
  signal type_cast_85_inst_ack_1 : boolean;
  signal type_cast_95_inst_req_0 : boolean;
  signal type_cast_95_inst_ack_0 : boolean;
  signal type_cast_95_inst_req_1 : boolean;
  signal type_cast_95_inst_ack_1 : boolean;
  signal type_cast_105_inst_req_0 : boolean;
  signal type_cast_105_inst_ack_0 : boolean;
  signal type_cast_105_inst_req_1 : boolean;
  signal type_cast_105_inst_ack_1 : boolean;
  signal type_cast_115_inst_req_0 : boolean;
  signal type_cast_115_inst_ack_0 : boolean;
  signal type_cast_115_inst_req_1 : boolean;
  signal type_cast_115_inst_ack_1 : boolean;
  signal type_cast_125_inst_req_0 : boolean;
  signal type_cast_125_inst_ack_0 : boolean;
  signal type_cast_125_inst_req_1 : boolean;
  signal type_cast_125_inst_ack_1 : boolean;
  signal type_cast_135_inst_req_0 : boolean;
  signal type_cast_135_inst_ack_0 : boolean;
  signal type_cast_135_inst_req_1 : boolean;
  signal type_cast_135_inst_ack_1 : boolean;
  signal type_cast_145_inst_req_0 : boolean;
  signal type_cast_145_inst_ack_0 : boolean;
  signal type_cast_145_inst_req_1 : boolean;
  signal type_cast_145_inst_ack_1 : boolean;
  signal type_cast_155_inst_req_0 : boolean;
  signal type_cast_155_inst_ack_0 : boolean;
  signal type_cast_155_inst_req_1 : boolean;
  signal type_cast_155_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_157_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_157_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_157_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_157_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_160_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_160_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_160_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_160_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_163_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_163_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_163_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_163_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_166_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_166_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_166_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_166_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_169_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_169_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_169_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_169_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_175_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_175_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_175_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_175_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_178_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_178_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_178_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_178_inst_ack_1 : boolean;
  signal if_stmt_192_branch_req_0 : boolean;
  signal if_stmt_192_branch_ack_1 : boolean;
  signal if_stmt_192_branch_ack_0 : boolean;
  signal phi_stmt_64_req_0 : boolean;
  signal type_cast_70_inst_req_0 : boolean;
  signal type_cast_70_inst_ack_0 : boolean;
  signal type_cast_70_inst_req_1 : boolean;
  signal type_cast_70_inst_ack_1 : boolean;
  signal phi_stmt_64_req_1 : boolean;
  signal phi_stmt_64_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_26: Block -- control-path 
    signal sendOutput_CP_26_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendOutput_CP_26_elements(0) <= sendOutput_CP_26_start;
    sendOutput_CP_26_symbol <= sendOutput_CP_26_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 branch_block_stmt_31/if_stmt_51_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_31/R_cmp68_52_place
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_31/$entry
      -- CP-element group 0: 	 branch_block_stmt_31/branch_block_stmt_31__entry__
      -- CP-element group 0: 	 branch_block_stmt_31/assign_stmt_41_to_assign_stmt_50__entry__
      -- CP-element group 0: 	 branch_block_stmt_31/assign_stmt_41_to_assign_stmt_50__exit__
      -- CP-element group 0: 	 branch_block_stmt_31/if_stmt_51__entry__
      -- CP-element group 0: 	 branch_block_stmt_31/assign_stmt_41_to_assign_stmt_50/$entry
      -- CP-element group 0: 	 branch_block_stmt_31/assign_stmt_41_to_assign_stmt_50/$exit
      -- CP-element group 0: 	 branch_block_stmt_31/if_stmt_51_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_31/if_stmt_51_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_31/if_stmt_51_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_31/if_stmt_51_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_31/if_stmt_51_else_link/$entry
      -- 
    branch_req_64_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_64_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => if_stmt_51_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	3 
    -- CP-element group 1: 	4 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_31/merge_stmt_57__exit__
      -- CP-element group 1: 	 branch_block_stmt_31/assign_stmt_61__entry__
      -- CP-element group 1: 	 branch_block_stmt_31/if_stmt_51_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_31/if_stmt_51_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_31/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_31/assign_stmt_61/$entry
      -- CP-element group 1: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_update_start_
      -- CP-element group 1: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_31/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_31/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_31/merge_stmt_57_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_31/merge_stmt_57_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_31/merge_stmt_57_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_31/merge_stmt_57_PhiAck/dummy
      -- 
    if_choice_transition_69_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_51_branch_ack_1, ack => sendOutput_CP_26_elements(1)); -- 
    rr_86_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_86_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(1), ack => type_cast_60_inst_req_0); -- 
    cr_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(1), ack => type_cast_60_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_31/if_stmt_51_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_31/if_stmt_51_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_31/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_31/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_31/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_73_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_51_branch_ack_0, ack => sendOutput_CP_26_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_Sample/ra
      -- 
    ra_87_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_60_inst_ack_0, ack => sendOutput_CP_26_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_31/assign_stmt_61__exit__
      -- CP-element group 4: 	 branch_block_stmt_31/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_31/assign_stmt_61/$exit
      -- CP-element group 4: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_31/assign_stmt_61/type_cast_60_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_31/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_31/bbx_xnph_forx_xbody_PhiReq/phi_stmt_64/$entry
      -- CP-element group 4: 	 branch_block_stmt_31/bbx_xnph_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/$entry
      -- 
    ca_92_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_60_inst_ack_1, ack => sendOutput_CP_26_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_final_index_sum_regn_Sample/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_76_index_offset_ack_0, ack => sendOutput_CP_26_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_request/req
      -- 
    ack_126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_76_index_offset_ack_1, ack => sendOutput_CP_26_elements(6)); -- 
    req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(6), ack => addr_of_77_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_request/$exit
      -- CP-element group 7: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_request/ack
      -- 
    ack_136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_77_final_reg_ack_0, ack => sendOutput_CP_26_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Sample/word_access_start/word_0/rr
      -- 
    ack_141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_77_final_reg_ack_1, ack => sendOutput_CP_26_elements(8)); -- 
    rr_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(8), ack => ptr_deref_81_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Sample/word_access_start/word_0/ra
      -- 
    ra_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_81_load_0_ack_0, ack => sendOutput_CP_26_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	21 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	25 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	17 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/ptr_deref_81_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/ptr_deref_81_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/ptr_deref_81_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/ptr_deref_81_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_Sample/rr
      -- 
    ca_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_81_load_0_ack_1, ack => sendOutput_CP_26_elements(10)); -- 
    rr_283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_145_inst_req_0); -- 
    rr_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_155_inst_req_0); -- 
    rr_213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_95_inst_req_0); -- 
    rr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_125_inst_req_0); -- 
    rr_241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_115_inst_req_0); -- 
    rr_199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_85_inst_req_0); -- 
    rr_269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_135_inst_req_0); -- 
    rr_227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_105_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_Sample/ra
      -- 
    ra_200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_0, ack => sendOutput_CP_26_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	47 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_Update/ca
      -- 
    ca_205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_1, ack => sendOutput_CP_26_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_Sample/ra
      -- 
    ra_214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_0, ack => sendOutput_CP_26_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	58 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	44 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_Update/ca
      -- 
    ca_219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_1, ack => sendOutput_CP_26_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_Sample/ra
      -- 
    ra_228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_105_inst_ack_0, ack => sendOutput_CP_26_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_Update/ca
      -- 
    ca_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_105_inst_ack_1, ack => sendOutput_CP_26_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_Sample/ra
      -- 
    ra_242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_115_inst_ack_0, ack => sendOutput_CP_26_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	58 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	38 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_Update/ca
      -- 
    ca_247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_115_inst_ack_1, ack => sendOutput_CP_26_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_Sample/ra
      -- 
    ra_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_125_inst_ack_0, ack => sendOutput_CP_26_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	58 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	35 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_Update/ca
      -- 
    ca_261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_125_inst_ack_1, ack => sendOutput_CP_26_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	10 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_Sample/ra
      -- 
    ra_270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_135_inst_ack_0, ack => sendOutput_CP_26_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	58 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	32 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_Update/ca
      -- 
    ca_275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_135_inst_ack_1, ack => sendOutput_CP_26_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_Sample/ra
      -- 
    ra_284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_0, ack => sendOutput_CP_26_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	58 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_Update/ca
      -- 
    ca_289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_1, ack => sendOutput_CP_26_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_Sample/ra
      -- 
    ra_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_0, ack => sendOutput_CP_26_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_Sample/req
      -- 
    ca_303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_1, ack => sendOutput_CP_26_elements(26)); -- 
    req_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(26), ack => WPIPE_zeropad_output_pipe_157_inst_req_0); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_update_start_
      -- CP-element group 27: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_Update/req
      -- 
    ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_157_inst_ack_0, ack => sendOutput_CP_26_elements(27)); -- 
    req_316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(27), ack => WPIPE_zeropad_output_pipe_157_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_157_Update/ack
      -- 
    ack_317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_157_inst_ack_1, ack => sendOutput_CP_26_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_Sample/req
      -- 
    req_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(29), ack => WPIPE_zeropad_output_pipe_160_inst_req_0); -- 
    sendOutput_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(24) & sendOutput_CP_26_elements(28);
      gj_sendOutput_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_update_start_
      -- CP-element group 30: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_Update/req
      -- 
    ack_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_160_inst_ack_0, ack => sendOutput_CP_26_elements(30)); -- 
    req_330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(30), ack => WPIPE_zeropad_output_pipe_160_inst_req_1); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_160_Update/ack
      -- 
    ack_331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_160_inst_ack_1, ack => sendOutput_CP_26_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	22 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_Sample/req
      -- 
    req_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(32), ack => WPIPE_zeropad_output_pipe_163_inst_req_0); -- 
    sendOutput_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(22) & sendOutput_CP_26_elements(31);
      gj_sendOutput_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_update_start_
      -- CP-element group 33: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_Update/req
      -- 
    ack_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_163_inst_ack_0, ack => sendOutput_CP_26_elements(33)); -- 
    req_344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(33), ack => WPIPE_zeropad_output_pipe_163_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_163_Update/ack
      -- 
    ack_345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_163_inst_ack_1, ack => sendOutput_CP_26_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	20 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_Sample/req
      -- 
    req_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(35), ack => WPIPE_zeropad_output_pipe_166_inst_req_0); -- 
    sendOutput_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(34) & sendOutput_CP_26_elements(20);
      gj_sendOutput_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_update_start_
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_Update/req
      -- 
    ack_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_166_inst_ack_0, ack => sendOutput_CP_26_elements(36)); -- 
    req_358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(36), ack => WPIPE_zeropad_output_pipe_166_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_166_Update/ack
      -- 
    ack_359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_166_inst_ack_1, ack => sendOutput_CP_26_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: 	18 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_Sample/req
      -- 
    req_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(38), ack => WPIPE_zeropad_output_pipe_169_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(37) & sendOutput_CP_26_elements(18);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_update_start_
      -- CP-element group 39: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_Update/req
      -- 
    ack_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_169_inst_ack_0, ack => sendOutput_CP_26_elements(39)); -- 
    req_372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(39), ack => WPIPE_zeropad_output_pipe_169_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_169_Update/ack
      -- 
    ack_373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_169_inst_ack_1, ack => sendOutput_CP_26_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: 	16 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_Sample/req
      -- 
    req_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(41), ack => WPIPE_zeropad_output_pipe_172_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(40) & sendOutput_CP_26_elements(16);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_update_start_
      -- CP-element group 42: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_Update/req
      -- 
    ack_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_172_inst_ack_0, ack => sendOutput_CP_26_elements(42)); -- 
    req_386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(42), ack => WPIPE_zeropad_output_pipe_172_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_172_Update/ack
      -- 
    ack_387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_172_inst_ack_1, ack => sendOutput_CP_26_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: 	14 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_Sample/req
      -- 
    req_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(44), ack => WPIPE_zeropad_output_pipe_175_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(43) & sendOutput_CP_26_elements(14);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_update_start_
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_Update/req
      -- 
    ack_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_175_inst_ack_0, ack => sendOutput_CP_26_elements(45)); -- 
    req_400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(45), ack => WPIPE_zeropad_output_pipe_175_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_175_Update/ack
      -- 
    ack_401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_175_inst_ack_1, ack => sendOutput_CP_26_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: 	12 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_Sample/req
      -- 
    req_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(47), ack => WPIPE_zeropad_output_pipe_178_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(46) & sendOutput_CP_26_elements(12);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_update_start_
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_Update/req
      -- 
    ack_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_178_inst_ack_0, ack => sendOutput_CP_26_elements(48)); -- 
    req_414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(48), ack => WPIPE_zeropad_output_pipe_178_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/WPIPE_zeropad_output_pipe_178_Update/ack
      -- 
    ack_415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_178_inst_ack_1, ack => sendOutput_CP_26_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	5 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191__exit__
      -- CP-element group 50: 	 branch_block_stmt_31/if_stmt_192__entry__
      -- CP-element group 50: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/$exit
      -- CP-element group 50: 	 branch_block_stmt_31/if_stmt_192_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/if_stmt_192_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/if_stmt_192_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_31/if_stmt_192_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_31/R_exitcond2_193_place
      -- CP-element group 50: 	 branch_block_stmt_31/if_stmt_192_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_31/if_stmt_192_else_link/$entry
      -- 
    branch_req_423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(50), ack => if_stmt_192_branch_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(49) & sendOutput_CP_26_elements(5);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_31/merge_stmt_198__exit__
      -- CP-element group 51: 	 branch_block_stmt_31/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_31/if_stmt_192_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_31/if_stmt_192_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_31/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_31/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_31/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_31/merge_stmt_198_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_31/merge_stmt_198_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_31/merge_stmt_198_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_31/merge_stmt_198_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_31/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_31/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_192_branch_ack_1, ack => sendOutput_CP_26_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_31/if_stmt_192_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_31/if_stmt_192_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_31/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/$entry
      -- CP-element group 52: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/$entry
      -- CP-element group 52: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/SplitProtocol/Update/cr
      -- 
    else_choice_transition_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_192_branch_ack_0, ack => sendOutput_CP_26_elements(52)); -- 
    rr_476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(52), ack => type_cast_70_inst_req_0); -- 
    cr_481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(52), ack => type_cast_70_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_31/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_31/bbx_xnph_forx_xbody_PhiReq/phi_stmt_64/$exit
      -- CP-element group 53: 	 branch_block_stmt_31/bbx_xnph_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_31/bbx_xnph_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_68_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_31/bbx_xnph_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_req
      -- 
    phi_stmt_64_req_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_64_req_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(53), ack => phi_stmt_64_req_0); -- 
    -- Element group sendOutput_CP_26_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendOutput_CP_26_elements(4), ack => sendOutput_CP_26_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/SplitProtocol/Sample/ra
      -- 
    ra_477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_70_inst_ack_0, ack => sendOutput_CP_26_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/SplitProtocol/Update/ca
      -- 
    ca_482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_70_inst_ack_1, ack => sendOutput_CP_26_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/$exit
      -- CP-element group 56: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/$exit
      -- CP-element group 56: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_sources/type_cast_70/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_31/forx_xbody_forx_xbody_PhiReq/phi_stmt_64/phi_stmt_64_req
      -- 
    phi_stmt_64_req_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_64_req_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(56), ack => phi_stmt_64_req_1); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(54) & sendOutput_CP_26_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	53 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_31/merge_stmt_63_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_31/merge_stmt_63_PhiAck/$entry
      -- 
    sendOutput_CP_26_elements(57) <= OrReduce(sendOutput_CP_26_elements(53) & sendOutput_CP_26_elements(56));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	22 
    -- CP-element group 58: 	24 
    -- CP-element group 58: 	26 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	12 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	10 
    -- CP-element group 58: 	14 
    -- CP-element group 58: 	20 
    -- CP-element group 58: 	18 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_31/merge_stmt_63__exit__
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191__entry__
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_update_start_
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/array_obj_ref_76_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/addr_of_77_complete/req
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_update_start_
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/ptr_deref_81_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_update_start_
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_85_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_update_start_
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_95_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_update_start_
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_105_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_update_start_
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_115_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_update_start_
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_125_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_update_start_
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_135_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_update_start_
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_145_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_update_start_
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_31/assign_stmt_78_to_assign_stmt_191/type_cast_155_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_31/merge_stmt_63_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_31/merge_stmt_63_PhiAck/phi_stmt_64_ack
      -- 
    phi_stmt_64_ack_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_64_ack_0, ack => sendOutput_CP_26_elements(58)); -- 
    cr_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => ptr_deref_81_load_0_req_1); -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => array_obj_ref_76_index_offset_req_0); -- 
    req_125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => array_obj_ref_76_index_offset_req_1); -- 
    req_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => addr_of_77_final_reg_req_1); -- 
    cr_204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_85_inst_req_1); -- 
    cr_218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_95_inst_req_1); -- 
    cr_232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_105_inst_req_1); -- 
    cr_246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_115_inst_req_1); -- 
    cr_260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_125_inst_req_1); -- 
    cr_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_135_inst_req_1); -- 
    cr_288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_145_inst_req_1); -- 
    cr_302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_155_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	51 
    -- CP-element group 59: 	2 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_31/$exit
      -- CP-element group 59: 	 branch_block_stmt_31/branch_block_stmt_31__exit__
      -- CP-element group 59: 	 branch_block_stmt_31/merge_stmt_200__exit__
      -- CP-element group 59: 	 branch_block_stmt_31/return__
      -- CP-element group 59: 	 branch_block_stmt_31/merge_stmt_202__exit__
      -- CP-element group 59: 	 branch_block_stmt_31/merge_stmt_200_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_31/merge_stmt_200_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_31/merge_stmt_200_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_31/merge_stmt_200_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_31/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_31/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_31/merge_stmt_202_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_31/merge_stmt_202_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_31/merge_stmt_202_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_31/merge_stmt_202_PhiAck/dummy
      -- 
    sendOutput_CP_26_elements(59) <= OrReduce(sendOutput_CP_26_elements(51) & sendOutput_CP_26_elements(2));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_39_wire : std_logic_vector(31 downto 0);
    signal R_indvar_75_resized : std_logic_vector(13 downto 0);
    signal R_indvar_75_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_76_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_76_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_76_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_76_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_76_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_76_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_78 : std_logic_vector(31 downto 0);
    signal cmp68_50 : std_logic_vector(0 downto 0);
    signal conv12_96 : std_logic_vector(7 downto 0);
    signal conv18_106 : std_logic_vector(7 downto 0);
    signal conv24_116 : std_logic_vector(7 downto 0);
    signal conv30_126 : std_logic_vector(7 downto 0);
    signal conv36_136 : std_logic_vector(7 downto 0);
    signal conv42_146 : std_logic_vector(7 downto 0);
    signal conv48_156 : std_logic_vector(7 downto 0);
    signal conv_86 : std_logic_vector(7 downto 0);
    signal exitcond2_191 : std_logic_vector(0 downto 0);
    signal indvar_64 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_186 : std_logic_vector(63 downto 0);
    signal ptr_deref_81_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_81_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_81_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_81_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_81_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_102 : std_logic_vector(63 downto 0);
    signal shr21_112 : std_logic_vector(63 downto 0);
    signal shr27_122 : std_logic_vector(63 downto 0);
    signal shr33_132 : std_logic_vector(63 downto 0);
    signal shr39_142 : std_logic_vector(63 downto 0);
    signal shr45_152 : std_logic_vector(63 downto 0);
    signal shr67_41 : std_logic_vector(31 downto 0);
    signal shr9_92 : std_logic_vector(63 downto 0);
    signal tmp1_61 : std_logic_vector(63 downto 0);
    signal tmp4_82 : std_logic_vector(63 downto 0);
    signal type_cast_100_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_110_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_120_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_130_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_140_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_150_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_184_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_35_wire : std_logic_vector(31 downto 0);
    signal type_cast_38_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_44_wire : std_logic_vector(31 downto 0);
    signal type_cast_47_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_68_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_70_wire : std_logic_vector(63 downto 0);
    signal type_cast_90_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_76_constant_part_of_offset <= "00000000000000";
    array_obj_ref_76_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_76_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_76_resized_base_address <= "00000000000000";
    ptr_deref_81_word_offset_0 <= "00000000000000";
    type_cast_100_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_110_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_120_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_130_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_140_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_150_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_184_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_38_wire_constant <= "00000000000000000000000000000010";
    type_cast_47_wire_constant <= "00000000000000000000000000000000";
    type_cast_68_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_90_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    phi_stmt_64: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_68_wire_constant & type_cast_70_wire;
      req <= phi_stmt_64_req_0 & phi_stmt_64_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_64",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_64_ack_0,
          idata => idata,
          odata => indvar_64,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_64
    addr_of_77_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_77_final_reg_req_0;
      addr_of_77_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_77_final_reg_req_1;
      addr_of_77_final_reg_ack_1<= rack(0);
      addr_of_77_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_77_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_76_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_78,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_105_inst_req_0;
      type_cast_105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_105_inst_req_1;
      type_cast_105_inst_ack_1<= rack(0);
      type_cast_105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_115_inst_req_0;
      type_cast_115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_115_inst_req_1;
      type_cast_115_inst_ack_1<= rack(0);
      type_cast_115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_115_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_116,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_125_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_125_inst_req_0;
      type_cast_125_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_125_inst_req_1;
      type_cast_125_inst_ack_1<= rack(0);
      type_cast_125_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_125_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_122,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_126,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_135_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_135_inst_req_0;
      type_cast_135_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_135_inst_req_1;
      type_cast_135_inst_ack_1<= rack(0);
      type_cast_135_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_135_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_136,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_145_inst_req_0;
      type_cast_145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_145_inst_req_1;
      type_cast_145_inst_ack_1<= rack(0);
      type_cast_145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_146,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_155_inst_req_0;
      type_cast_155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_155_inst_req_1;
      type_cast_155_inst_ack_1<= rack(0);
      type_cast_155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_152,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_156,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_35_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := size_buffer(31 downto 0);
      type_cast_35_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_40_inst
    process(ASHR_i32_i32_39_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_39_wire(31 downto 0);
      shr67_41 <= tmp_var; -- 
    end process;
    -- interlock type_cast_44_inst
    process(shr67_41) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := shr67_41(31 downto 0);
      type_cast_44_wire <= tmp_var; -- 
    end process;
    type_cast_60_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_60_inst_req_0;
      type_cast_60_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_60_inst_req_1;
      type_cast_60_inst_ack_1<= rack(0);
      type_cast_60_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_60_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr67_41,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_61,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_70_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_70_inst_req_0;
      type_cast_70_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_70_inst_req_1;
      type_cast_70_inst_ack_1<= rack(0);
      type_cast_70_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_70_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_70_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_85_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_85_inst_req_0;
      type_cast_85_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_85_inst_req_1;
      type_cast_85_inst_ack_1<= rack(0);
      type_cast_85_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_85_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_82,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_86,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_95_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_95_inst_req_0;
      type_cast_95_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_95_inst_req_1;
      type_cast_95_inst_ack_1<= rack(0);
      type_cast_95_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_95_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_92,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_96,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_76_index_1_rename
    process(R_indvar_75_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_75_resized;
      ov(13 downto 0) := iv;
      R_indvar_75_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_76_index_1_resize
    process(indvar_64) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_64;
      ov := iv(13 downto 0);
      R_indvar_75_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_76_root_address_inst
    process(array_obj_ref_76_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_76_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_76_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_81_addr_0
    process(ptr_deref_81_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_81_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_81_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_81_base_resize
    process(arrayidx_78) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_78;
      ov := iv(13 downto 0);
      ptr_deref_81_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_81_gather_scatter
    process(ptr_deref_81_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_81_data_0;
      ov(63 downto 0) := iv;
      tmp4_82 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_81_root_address_inst
    process(ptr_deref_81_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_81_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_81_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_192_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_191;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_192_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_192_branch_req_0,
          ack0 => if_stmt_192_branch_ack_0,
          ack1 => if_stmt_192_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_51_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp68_50;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_51_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_51_branch_req_0,
          ack0 => if_stmt_51_branch_ack_0,
          ack1 => if_stmt_51_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_185_inst
    process(indvar_64) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_64, type_cast_184_wire_constant, tmp_var);
      indvarx_xnext_186 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_39_inst
    process(type_cast_35_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_35_wire, type_cast_38_wire_constant, tmp_var);
      ASHR_i32_i32_39_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_190_inst
    process(indvarx_xnext_186, tmp1_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_186, tmp1_61, tmp_var);
      exitcond2_191 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_101_inst
    process(tmp4_82) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_82, type_cast_100_wire_constant, tmp_var);
      shr15_102 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_111_inst
    process(tmp4_82) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_82, type_cast_110_wire_constant, tmp_var);
      shr21_112 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_121_inst
    process(tmp4_82) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_82, type_cast_120_wire_constant, tmp_var);
      shr27_122 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_131_inst
    process(tmp4_82) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_82, type_cast_130_wire_constant, tmp_var);
      shr33_132 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_141_inst
    process(tmp4_82) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_82, type_cast_140_wire_constant, tmp_var);
      shr39_142 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_151_inst
    process(tmp4_82) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_82, type_cast_150_wire_constant, tmp_var);
      shr45_152 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_91_inst
    process(tmp4_82) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_82, type_cast_90_wire_constant, tmp_var);
      shr9_92 <= tmp_var; --
    end process;
    -- binary operator SGT_i32_u1_48_inst
    process(type_cast_44_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(type_cast_44_wire, type_cast_47_wire_constant, tmp_var);
      cmp68_50 <= tmp_var; --
    end process;
    -- shared split operator group (11) : array_obj_ref_76_index_offset 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_75_scaled;
      array_obj_ref_76_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_76_index_offset_req_0;
      array_obj_ref_76_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_76_index_offset_req_1;
      array_obj_ref_76_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_11_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared load operator group (0) : ptr_deref_81_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_81_load_0_req_0;
      ptr_deref_81_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_81_load_0_req_1;
      ptr_deref_81_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_81_word_address_0;
      ptr_deref_81_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_157_inst WPIPE_zeropad_output_pipe_160_inst WPIPE_zeropad_output_pipe_163_inst WPIPE_zeropad_output_pipe_166_inst WPIPE_zeropad_output_pipe_169_inst WPIPE_zeropad_output_pipe_172_inst WPIPE_zeropad_output_pipe_175_inst WPIPE_zeropad_output_pipe_178_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_157_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_160_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_163_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_166_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_169_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_172_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_175_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_178_inst_req_0;
      WPIPE_zeropad_output_pipe_157_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_160_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_163_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_166_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_169_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_172_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_175_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_178_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_157_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_160_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_163_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_166_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_169_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_172_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_175_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_178_inst_req_1;
      WPIPE_zeropad_output_pipe_157_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_160_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_163_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_166_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_169_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_172_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_175_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_178_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv48_156 & conv42_146 & conv36_136 & conv30_126 & conv24_116 & conv18_106 & conv12_96 & conv_86;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_520_start: Boolean;
  signal timer_CP_520_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_208_load_0_req_0 : boolean;
  signal LOAD_count_208_load_0_ack_0 : boolean;
  signal LOAD_count_208_load_0_req_1 : boolean;
  signal LOAD_count_208_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_520_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_520_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_520_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_520_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_520: Block -- control-path 
    signal timer_CP_520_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_520_elements(0) <= timer_CP_520_start;
    timer_CP_520_symbol <= timer_CP_520_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_209/$entry
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_sample_start_
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_update_start_
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_Update/$entry
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_209/LOAD_count_208_Update/word_access_complete/word_0/cr
      -- 
    cr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_520_elements(0), ack => LOAD_count_208_load_0_req_1); -- 
    rr_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_520_elements(0), ack => LOAD_count_208_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_209/LOAD_count_208_sample_completed_
      -- CP-element group 1: 	 assign_stmt_209/LOAD_count_208_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_209/LOAD_count_208_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_209/LOAD_count_208_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_209/LOAD_count_208_Sample/word_access_start/word_0/ra
      -- 
    ra_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_208_load_0_ack_0, ack => timer_CP_520_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_209/$exit
      -- CP-element group 2: 	 assign_stmt_209/LOAD_count_208_update_completed_
      -- CP-element group 2: 	 assign_stmt_209/LOAD_count_208_Update/$exit
      -- CP-element group 2: 	 assign_stmt_209/LOAD_count_208_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_209/LOAD_count_208_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_209/LOAD_count_208_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_209/LOAD_count_208_Update/LOAD_count_208_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_209/LOAD_count_208_Update/LOAD_count_208_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_209/LOAD_count_208_Update/LOAD_count_208_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_209/LOAD_count_208_Update/LOAD_count_208_Merge/merge_ack
      -- 
    ca_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_208_load_0_ack_1, ack => timer_CP_520_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_208_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_208_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_208_word_address_0 <= "0";
    -- equivalence LOAD_count_208_gather_scatter
    process(LOAD_count_208_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_208_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_208_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_208_load_0_req_0;
      LOAD_count_208_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_208_load_0_req_1;
      LOAD_count_208_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_208_word_address_0;
      LOAD_count_208_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block1_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block3_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block1_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block0_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block3_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    Block2_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_data : out  std_logic_vector(31 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D;
architecture zeropad3D_arch of zeropad3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_CP_676_start: Boolean;
  signal zeropad3D_CP_676_symbol: Boolean;
  -- volatile/operator module components. 
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_zeropad_input_pipe_248_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_257_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_633_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_566_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_554_inst_req_0 : boolean;
  signal type_cast_306_inst_req_1 : boolean;
  signal type_cast_306_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_566_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_248_inst_ack_0 : boolean;
  signal WPIPE_Block3_starting_587_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_563_inst_req_1 : boolean;
  signal RPIPE_Block0_complete_609_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_584_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_242_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_239_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_566_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_242_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_236_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_563_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_563_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_239_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_587_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_584_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_236_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_236_inst_req_1 : boolean;
  signal WPIPE_Block1_starting_551_inst_ack_0 : boolean;
  signal type_cast_261_inst_ack_0 : boolean;
  signal RPIPE_Block0_complete_609_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_569_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_593_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_569_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_572_inst_ack_0 : boolean;
  signal WPIPE_Block3_starting_587_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_554_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_233_inst_ack_0 : boolean;
  signal type_cast_261_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_233_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_602_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_593_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_560_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_602_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_239_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_593_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_551_inst_req_0 : boolean;
  signal type_cast_643_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_236_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_245_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_245_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_569_inst_req_0 : boolean;
  signal WPIPE_Block2_starting_572_inst_req_0 : boolean;
  signal RPIPE_Block2_complete_615_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_563_inst_ack_0 : boolean;
  signal if_stmt_293_branch_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_633_inst_req_1 : boolean;
  signal type_cast_643_inst_req_0 : boolean;
  signal type_cast_306_inst_ack_0 : boolean;
  signal type_cast_265_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_581_inst_req_1 : boolean;
  signal RPIPE_Block2_complete_615_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_233_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_593_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_245_inst_ack_0 : boolean;
  signal type_cast_626_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_596_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_566_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_239_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_584_inst_req_1 : boolean;
  signal type_cast_626_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_554_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_245_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_233_inst_ack_1 : boolean;
  signal if_stmt_293_branch_req_0 : boolean;
  signal type_cast_269_inst_ack_1 : boolean;
  signal type_cast_269_inst_req_1 : boolean;
  signal type_cast_269_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_0 : boolean;
  signal type_cast_265_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_254_inst_ack_1 : boolean;
  signal type_cast_261_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_254_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_254_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_254_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_602_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_602_inst_ack_0 : boolean;
  signal type_cast_265_inst_ack_0 : boolean;
  signal RPIPE_Block0_complete_609_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_257_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_560_inst_ack_1 : boolean;
  signal call_stmt_660_call_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_251_inst_ack_0 : boolean;
  signal if_stmt_293_branch_ack_1 : boolean;
  signal type_cast_643_inst_ack_0 : boolean;
  signal RPIPE_Block0_complete_609_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_251_inst_req_0 : boolean;
  signal WPIPE_Block2_starting_584_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_248_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_248_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_596_inst_req_0 : boolean;
  signal type_cast_265_inst_req_1 : boolean;
  signal WPIPE_Block1_starting_554_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_257_inst_ack_1 : boolean;
  signal type_cast_261_inst_ack_1 : boolean;
  signal type_cast_626_inst_ack_0 : boolean;
  signal WPIPE_Block3_starting_590_inst_ack_1 : boolean;
  signal type_cast_315_inst_req_1 : boolean;
  signal type_cast_315_inst_ack_1 : boolean;
  signal type_cast_315_inst_req_0 : boolean;
  signal type_cast_315_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_242_inst_ack_0 : boolean;
  signal call_stmt_622_call_ack_1 : boolean;
  signal WPIPE_Block2_starting_581_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_569_inst_ack_0 : boolean;
  signal WPIPE_Block3_starting_590_inst_req_1 : boolean;
  signal type_cast_302_inst_req_0 : boolean;
  signal type_cast_302_inst_ack_0 : boolean;
  signal type_cast_626_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_242_inst_req_0 : boolean;
  signal type_cast_647_inst_req_1 : boolean;
  signal phi_stmt_343_req_0 : boolean;
  signal type_cast_647_inst_ack_1 : boolean;
  signal type_cast_302_inst_ack_1 : boolean;
  signal type_cast_302_inst_req_1 : boolean;
  signal type_cast_306_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_251_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_257_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_251_inst_req_1 : boolean;
  signal RPIPE_Block2_complete_615_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_587_inst_req_1 : boolean;
  signal WPIPE_Block2_starting_581_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_581_inst_req_0 : boolean;
  signal type_cast_647_inst_ack_0 : boolean;
  signal WPIPE_Block3_starting_590_inst_ack_0 : boolean;
  signal call_stmt_622_call_req_1 : boolean;
  signal RPIPE_Block1_complete_612_inst_ack_1 : boolean;
  signal array_obj_ref_355_index_offset_req_0 : boolean;
  signal array_obj_ref_355_index_offset_ack_0 : boolean;
  signal array_obj_ref_355_index_offset_req_1 : boolean;
  signal array_obj_ref_355_index_offset_ack_1 : boolean;
  signal RPIPE_Block2_complete_615_inst_req_1 : boolean;
  signal call_stmt_660_call_ack_0 : boolean;
  signal WPIPE_Block1_starting_560_inst_ack_0 : boolean;
  signal addr_of_356_final_reg_req_0 : boolean;
  signal addr_of_356_final_reg_ack_0 : boolean;
  signal addr_of_356_final_reg_req_1 : boolean;
  signal addr_of_356_final_reg_ack_1 : boolean;
  signal RPIPE_Block1_complete_612_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_590_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_359_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_359_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_560_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_359_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_359_inst_ack_1 : boolean;
  signal type_cast_647_inst_req_0 : boolean;
  signal call_stmt_622_call_ack_0 : boolean;
  signal type_cast_363_inst_req_0 : boolean;
  signal type_cast_363_inst_ack_0 : boolean;
  signal type_cast_363_inst_req_1 : boolean;
  signal type_cast_363_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_372_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_372_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_372_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_372_inst_ack_1 : boolean;
  signal call_stmt_622_call_req_0 : boolean;
  signal type_cast_376_inst_req_0 : boolean;
  signal type_cast_376_inst_ack_0 : boolean;
  signal type_cast_376_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_599_inst_ack_1 : boolean;
  signal type_cast_376_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_633_inst_ack_0 : boolean;
  signal RPIPE_Block1_complete_612_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_390_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_390_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_390_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_599_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_390_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_578_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_578_inst_req_1 : boolean;
  signal type_cast_394_inst_req_0 : boolean;
  signal type_cast_394_inst_ack_0 : boolean;
  signal type_cast_394_inst_req_1 : boolean;
  signal type_cast_394_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_633_inst_req_0 : boolean;
  signal RPIPE_Block1_complete_612_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_408_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_408_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_408_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_408_inst_ack_1 : boolean;
  signal type_cast_412_inst_req_0 : boolean;
  signal type_cast_412_inst_ack_0 : boolean;
  signal type_cast_412_inst_req_1 : boolean;
  signal WPIPE_Block1_starting_548_inst_ack_1 : boolean;
  signal type_cast_412_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_599_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_426_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_426_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_426_inst_req_1 : boolean;
  signal WPIPE_Block3_starting_599_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_426_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_578_inst_ack_0 : boolean;
  signal WPIPE_Block2_starting_578_inst_req_0 : boolean;
  signal type_cast_430_inst_req_0 : boolean;
  signal type_cast_430_inst_ack_0 : boolean;
  signal type_cast_430_inst_req_1 : boolean;
  signal type_cast_430_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_444_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_444_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_444_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_444_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_605_inst_ack_1 : boolean;
  signal type_cast_448_inst_req_0 : boolean;
  signal type_cast_448_inst_ack_0 : boolean;
  signal RPIPE_Block3_complete_618_inst_ack_1 : boolean;
  signal type_cast_448_inst_req_1 : boolean;
  signal type_cast_448_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_605_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_462_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_462_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_462_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_462_inst_ack_1 : boolean;
  signal call_stmt_660_call_ack_1 : boolean;
  signal RPIPE_Block3_complete_618_inst_req_1 : boolean;
  signal type_cast_466_inst_req_0 : boolean;
  signal type_cast_466_inst_ack_0 : boolean;
  signal type_cast_466_inst_req_1 : boolean;
  signal type_cast_466_inst_ack_1 : boolean;
  signal type_cast_639_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_480_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_480_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_557_inst_ack_1 : boolean;
  signal type_cast_639_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_480_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_480_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_605_inst_ack_0 : boolean;
  signal type_cast_484_inst_req_0 : boolean;
  signal type_cast_484_inst_ack_0 : boolean;
  signal type_cast_484_inst_req_1 : boolean;
  signal type_cast_484_inst_ack_1 : boolean;
  signal WPIPE_Block3_starting_605_inst_req_0 : boolean;
  signal WPIPE_Block2_starting_575_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_575_inst_req_1 : boolean;
  signal ptr_deref_492_store_0_req_0 : boolean;
  signal ptr_deref_492_store_0_ack_0 : boolean;
  signal ptr_deref_492_store_0_req_1 : boolean;
  signal WPIPE_Block2_starting_575_inst_ack_0 : boolean;
  signal ptr_deref_492_store_0_ack_1 : boolean;
  signal WPIPE_Block2_starting_575_inst_req_0 : boolean;
  signal call_stmt_660_call_req_0 : boolean;
  signal RPIPE_Block3_complete_618_inst_ack_0 : boolean;
  signal if_stmt_506_branch_req_0 : boolean;
  signal WPIPE_Block1_starting_551_inst_ack_1 : boolean;
  signal if_stmt_506_branch_ack_1 : boolean;
  signal WPIPE_Block1_starting_551_inst_req_1 : boolean;
  signal if_stmt_506_branch_ack_0 : boolean;
  signal WPIPE_Block1_starting_548_inst_req_1 : boolean;
  signal type_cast_639_inst_ack_0 : boolean;
  signal call_stmt_517_call_req_0 : boolean;
  signal call_stmt_517_call_ack_0 : boolean;
  signal RPIPE_Block3_complete_618_inst_req_0 : boolean;
  signal call_stmt_517_call_req_1 : boolean;
  signal call_stmt_517_call_ack_1 : boolean;
  signal type_cast_522_inst_req_0 : boolean;
  signal type_cast_522_inst_ack_0 : boolean;
  signal type_cast_522_inst_req_1 : boolean;
  signal type_cast_522_inst_ack_1 : boolean;
  signal type_cast_639_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_524_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_596_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_524_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_524_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_524_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_557_inst_req_1 : boolean;
  signal type_cast_643_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_527_inst_req_0 : boolean;
  signal WPIPE_Block3_starting_596_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_527_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_527_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_527_inst_ack_1 : boolean;
  signal WPIPE_Block2_starting_572_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_530_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_530_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_557_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_530_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_530_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_557_inst_req_0 : boolean;
  signal WPIPE_Block2_starting_572_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_533_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_533_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_533_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_533_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_536_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_536_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_536_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_536_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_539_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_539_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_539_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_539_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_542_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_542_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_542_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_542_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_545_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_545_inst_ack_0 : boolean;
  signal WPIPE_Block1_starting_545_inst_req_1 : boolean;
  signal WPIPE_Block1_starting_545_inst_ack_1 : boolean;
  signal WPIPE_Block1_starting_548_inst_req_0 : boolean;
  signal WPIPE_Block1_starting_548_inst_ack_0 : boolean;
  signal type_cast_349_inst_req_0 : boolean;
  signal type_cast_349_inst_ack_0 : boolean;
  signal type_cast_349_inst_req_1 : boolean;
  signal type_cast_349_inst_ack_1 : boolean;
  signal phi_stmt_343_req_1 : boolean;
  signal phi_stmt_343_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_CP_676_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_676_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_CP_676_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_676_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_CP_676: Block -- control-path 
    signal zeropad3D_CP_676_elements: BooleanArray(167 downto 0);
    -- 
  begin -- 
    zeropad3D_CP_676_elements(0) <= zeropad3D_CP_676_start;
    zeropad3D_CP_676_symbol <= zeropad3D_CP_676_elements(160);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	22 
    -- CP-element group 0: 	24 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/$entry
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_update_start_
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292__entry__
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_231/branch_block_stmt_231__entry__
      -- CP-element group 0: 	 branch_block_stmt_231/$entry
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_update_start_
      -- CP-element group 0: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_update_start_
      -- 
    rr_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => RPIPE_zeropad_input_pipe_233_inst_req_0); -- 
    cr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_269_inst_req_1); -- 
    cr_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_261_inst_req_1); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_265_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_update_start_
      -- CP-element group 1: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_Sample/$exit
      -- 
    ra_721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_233_inst_ack_0, ack => zeropad3D_CP_676_elements(1)); -- 
    cr_725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(1), ack => RPIPE_zeropad_input_pipe_233_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_233_Update/ca
      -- 
    ca_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_233_inst_ack_1, ack => zeropad3D_CP_676_elements(2)); -- 
    rr_734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(2), ack => RPIPE_zeropad_input_pipe_236_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_update_start_
      -- CP-element group 3: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_sample_completed_
      -- 
    ra_735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_236_inst_ack_0, ack => zeropad3D_CP_676_elements(3)); -- 
    cr_739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(3), ack => RPIPE_zeropad_input_pipe_236_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_236_update_completed_
      -- 
    ca_740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_236_inst_ack_1, ack => zeropad3D_CP_676_elements(4)); -- 
    rr_748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(4), ack => RPIPE_zeropad_input_pipe_239_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_update_start_
      -- CP-element group 5: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_Update/$entry
      -- 
    ra_749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_239_inst_ack_0, ack => zeropad3D_CP_676_elements(5)); -- 
    cr_753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(5), ack => RPIPE_zeropad_input_pipe_239_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	19 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_239_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_Sample/$entry
      -- 
    ca_754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_239_inst_ack_1, ack => zeropad3D_CP_676_elements(6)); -- 
    rr_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => RPIPE_zeropad_input_pipe_242_inst_req_0); -- 
    rr_846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => type_cast_261_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_update_start_
      -- CP-element group 7: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_Sample/$exit
      -- 
    ra_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_242_inst_ack_0, ack => zeropad3D_CP_676_elements(7)); -- 
    cr_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(7), ack => RPIPE_zeropad_input_pipe_242_inst_req_1); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_242_update_completed_
      -- 
    ca_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_242_inst_ack_1, ack => zeropad3D_CP_676_elements(8)); -- 
    rr_776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => RPIPE_zeropad_input_pipe_245_inst_req_0); -- 
    rr_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => type_cast_265_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_update_start_
      -- CP-element group 9: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_Sample/$exit
      -- 
    ra_777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_245_inst_ack_0, ack => zeropad3D_CP_676_elements(9)); -- 
    cr_781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(9), ack => RPIPE_zeropad_input_pipe_245_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	23 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_245_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_Sample/$entry
      -- 
    ca_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_245_inst_ack_1, ack => zeropad3D_CP_676_elements(10)); -- 
    rr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(10), ack => RPIPE_zeropad_input_pipe_248_inst_req_0); -- 
    rr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(10), ack => type_cast_269_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_update_start_
      -- CP-element group 11: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_Update/$entry
      -- 
    ra_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_248_inst_ack_0, ack => zeropad3D_CP_676_elements(11)); -- 
    cr_795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(11), ack => RPIPE_zeropad_input_pipe_248_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_248_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_sample_start_
      -- 
    ca_796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_248_inst_ack_1, ack => zeropad3D_CP_676_elements(12)); -- 
    rr_804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(12), ack => RPIPE_zeropad_input_pipe_251_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_update_start_
      -- CP-element group 13: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_Update/cr
      -- 
    ra_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_251_inst_ack_0, ack => zeropad3D_CP_676_elements(13)); -- 
    cr_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(13), ack => RPIPE_zeropad_input_pipe_251_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_251_Update/ca
      -- 
    ca_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_251_inst_ack_1, ack => zeropad3D_CP_676_elements(14)); -- 
    rr_818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(14), ack => RPIPE_zeropad_input_pipe_254_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_update_start_
      -- CP-element group 15: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_sample_completed_
      -- 
    ra_819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_254_inst_ack_0, ack => zeropad3D_CP_676_elements(15)); -- 
    cr_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(15), ack => RPIPE_zeropad_input_pipe_254_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_254_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_Sample/$entry
      -- 
    ca_824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_254_inst_ack_1, ack => zeropad3D_CP_676_elements(16)); -- 
    rr_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(16), ack => RPIPE_zeropad_input_pipe_257_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_update_start_
      -- CP-element group 17: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_Update/cr
      -- 
    ra_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_257_inst_ack_0, ack => zeropad3D_CP_676_elements(17)); -- 
    cr_837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(17), ack => RPIPE_zeropad_input_pipe_257_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	25 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/RPIPE_zeropad_input_pipe_257_update_completed_
      -- 
    ca_838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_257_inst_ack_1, ack => zeropad3D_CP_676_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	6 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_sample_completed_
      -- 
    ra_847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_0, ack => zeropad3D_CP_676_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	25 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_261_Update/ca
      -- 
    ca_852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_1, ack => zeropad3D_CP_676_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_Sample/$exit
      -- 
    ra_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_0, ack => zeropad3D_CP_676_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	0 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_265_update_completed_
      -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_1, ack => zeropad3D_CP_676_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_Sample/$exit
      -- 
    ra_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_0, ack => zeropad3D_CP_676_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/type_cast_269_update_completed_
      -- 
    ca_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_1, ack => zeropad3D_CP_676_elements(24)); -- 
    -- CP-element group 25:  branch  join  transition  place  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: 	20 
    -- CP-element group 25: 	22 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (10) 
      -- CP-element group 25: 	 branch_block_stmt_231/if_stmt_293_if_link/$entry
      -- CP-element group 25: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292/$exit
      -- CP-element group 25: 	 branch_block_stmt_231/if_stmt_293__entry__
      -- CP-element group 25: 	 branch_block_stmt_231/assign_stmt_234_to_assign_stmt_292__exit__
      -- CP-element group 25: 	 branch_block_stmt_231/if_stmt_293_dead_link/$entry
      -- CP-element group 25: 	 branch_block_stmt_231/if_stmt_293_eval_test/branch_req
      -- CP-element group 25: 	 branch_block_stmt_231/if_stmt_293_eval_test/$entry
      -- CP-element group 25: 	 branch_block_stmt_231/if_stmt_293_eval_test/$exit
      -- CP-element group 25: 	 branch_block_stmt_231/R_cmp126_294_place
      -- CP-element group 25: 	 branch_block_stmt_231/if_stmt_293_else_link/$entry
      -- 
    branch_req_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(25), ack => if_stmt_293_branch_req_0); -- 
    zeropad3D_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(18) & zeropad3D_CP_676_elements(20) & zeropad3D_CP_676_elements(22) & zeropad3D_CP_676_elements(24);
      gj_zeropad3D_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  place  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	167 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_231/if_stmt_293_if_link/$exit
      -- CP-element group 26: 	 branch_block_stmt_231/if_stmt_293_if_link/if_choice_transition
      -- CP-element group 26: 	 branch_block_stmt_231/entry_forx_xend
      -- CP-element group 26: 	 branch_block_stmt_231/entry_forx_xend_PhiReq/$entry
      -- CP-element group 26: 	 branch_block_stmt_231/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_293_branch_ack_1, ack => zeropad3D_CP_676_elements(26)); -- 
    -- CP-element group 27:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	29 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	31 
    -- CP-element group 27: 	32 
    -- CP-element group 27: 	33 
    -- CP-element group 27:  members (30) 
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340__entry__
      -- CP-element group 27: 	 branch_block_stmt_231/merge_stmt_299__exit__
      -- CP-element group 27: 	 branch_block_stmt_231/if_stmt_293_else_link/else_choice_transition
      -- CP-element group 27: 	 branch_block_stmt_231/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_update_start_
      -- CP-element group 27: 	 branch_block_stmt_231/entry_bbx_xnph
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_update_start_
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_231/if_stmt_293_else_link/$exit
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/$entry
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_update_start_
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_231/merge_stmt_299_PhiAck/dummy
      -- CP-element group 27: 	 branch_block_stmt_231/merge_stmt_299_PhiAck/$exit
      -- CP-element group 27: 	 branch_block_stmt_231/merge_stmt_299_PhiAck/$entry
      -- CP-element group 27: 	 branch_block_stmt_231/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 27: 	 branch_block_stmt_231/merge_stmt_299_PhiReqMerge
      -- 
    else_choice_transition_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_293_branch_ack_0, ack => zeropad3D_CP_676_elements(27)); -- 
    cr_929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_306_inst_req_1); -- 
    cr_943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_315_inst_req_1); -- 
    rr_938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_315_inst_req_0); -- 
    rr_910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_302_inst_req_0); -- 
    cr_915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_302_inst_req_1); -- 
    rr_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => type_cast_306_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_Sample/ra
      -- 
    ra_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_0, ack => zeropad3D_CP_676_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_302_Update/$exit
      -- 
    ca_916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_1, ack => zeropad3D_CP_676_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_Sample/$exit
      -- 
    ra_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_306_inst_ack_0, ack => zeropad3D_CP_676_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	27 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_306_update_completed_
      -- 
    ca_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_306_inst_ack_1, ack => zeropad3D_CP_676_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	27 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_Sample/ra
      -- 
    ra_939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_315_inst_ack_0, ack => zeropad3D_CP_676_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	27 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/type_cast_315_update_completed_
      -- 
    ca_944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_315_inst_ack_1, ack => zeropad3D_CP_676_elements(33)); -- 
    -- CP-element group 34:  join  transition  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	161 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_231/bbx_xnph_forx_xbody
      -- CP-element group 34: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340__exit__
      -- CP-element group 34: 	 branch_block_stmt_231/assign_stmt_303_to_assign_stmt_340/$exit
      -- CP-element group 34: 	 branch_block_stmt_231/bbx_xnph_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_231/bbx_xnph_forx_xbody_PhiReq/phi_stmt_343/$entry
      -- CP-element group 34: 	 branch_block_stmt_231/bbx_xnph_forx_xbody_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(29) & zeropad3D_CP_676_elements(31) & zeropad3D_CP_676_elements(33);
      gj_zeropad3D_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	166 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	74 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_final_index_sum_regn_sample_complete
      -- CP-element group 35: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_final_index_sum_regn_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_final_index_sum_regn_Sample/ack
      -- 
    ack_973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_355_index_offset_ack_0, ack => zeropad3D_CP_676_elements(35)); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	166 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (11) 
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_root_address_calculated
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_offset_calculated
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_final_index_sum_regn_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_final_index_sum_regn_Update/ack
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_base_plus_offset/$entry
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_base_plus_offset/$exit
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_base_plus_offset/sum_rename_req
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_base_plus_offset/sum_rename_ack
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_request/$entry
      -- CP-element group 36: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_request/req
      -- 
    ack_978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_355_index_offset_ack_1, ack => zeropad3D_CP_676_elements(36)); -- 
    req_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(36), ack => addr_of_356_final_reg_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_request/$exit
      -- CP-element group 37: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_request/ack
      -- 
    ack_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_356_final_reg_ack_0, ack => zeropad3D_CP_676_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	166 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	71 
    -- CP-element group 38:  members (19) 
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_complete/$exit
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_complete/ack
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_base_address_calculated
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_word_address_calculated
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_root_address_calculated
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_base_address_resized
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_base_addr_resize/$entry
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_base_addr_resize/$exit
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_base_addr_resize/base_resize_req
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_base_addr_resize/base_resize_ack
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_base_plus_offset/$entry
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_base_plus_offset/$exit
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_base_plus_offset/sum_rename_req
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_base_plus_offset/sum_rename_ack
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_word_addrgen/$entry
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_word_addrgen/$exit
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_word_addrgen/root_register_req
      -- CP-element group 38: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_word_addrgen/root_register_ack
      -- 
    ack_993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_356_final_reg_ack_1, ack => zeropad3D_CP_676_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	166 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_update_start_
      -- CP-element group 39: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_Update/cr
      -- 
    ra_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_359_inst_ack_0, ack => zeropad3D_CP_676_elements(39)); -- 
    cr_1006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(39), ack => RPIPE_zeropad_input_pipe_359_inst_req_1); -- 
    -- CP-element group 40:  fork  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_Sample/rr
      -- CP-element group 40: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_Sample/rr
      -- 
    ca_1007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_359_inst_ack_1, ack => zeropad3D_CP_676_elements(40)); -- 
    rr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(40), ack => type_cast_363_inst_req_0); -- 
    rr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(40), ack => RPIPE_zeropad_input_pipe_372_inst_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_Sample/ra
      -- 
    ra_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_363_inst_ack_0, ack => zeropad3D_CP_676_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	166 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	71 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_Update/ca
      -- 
    ca_1021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_363_inst_ack_1, ack => zeropad3D_CP_676_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	40 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_update_start_
      -- CP-element group 43: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_Update/cr
      -- 
    ra_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_372_inst_ack_0, ack => zeropad3D_CP_676_elements(43)); -- 
    cr_1034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(43), ack => RPIPE_zeropad_input_pipe_372_inst_req_1); -- 
    -- CP-element group 44:  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_372_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_Sample/rr
      -- CP-element group 44: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_Sample/rr
      -- 
    ca_1035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_372_inst_ack_1, ack => zeropad3D_CP_676_elements(44)); -- 
    rr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(44), ack => type_cast_376_inst_req_0); -- 
    rr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(44), ack => RPIPE_zeropad_input_pipe_390_inst_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_Sample/ra
      -- 
    ra_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_376_inst_ack_0, ack => zeropad3D_CP_676_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	166 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	71 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_Update/ca
      -- 
    ca_1049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_376_inst_ack_1, ack => zeropad3D_CP_676_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_update_start_
      -- CP-element group 47: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_Update/cr
      -- 
    ra_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_390_inst_ack_0, ack => zeropad3D_CP_676_elements(47)); -- 
    cr_1062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(47), ack => RPIPE_zeropad_input_pipe_390_inst_req_1); -- 
    -- CP-element group 48:  fork  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: 	51 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_390_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_Sample/rr
      -- CP-element group 48: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_Sample/rr
      -- 
    ca_1063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_390_inst_ack_1, ack => zeropad3D_CP_676_elements(48)); -- 
    rr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(48), ack => type_cast_394_inst_req_0); -- 
    rr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(48), ack => RPIPE_zeropad_input_pipe_408_inst_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_Sample/ra
      -- 
    ra_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_394_inst_ack_0, ack => zeropad3D_CP_676_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	166 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	71 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_Update/ca
      -- 
    ca_1077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_394_inst_ack_1, ack => zeropad3D_CP_676_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	48 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_update_start_
      -- CP-element group 51: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_Update/cr
      -- 
    ra_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_408_inst_ack_0, ack => zeropad3D_CP_676_elements(51)); -- 
    cr_1090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(51), ack => RPIPE_zeropad_input_pipe_408_inst_req_1); -- 
    -- CP-element group 52:  fork  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (9) 
      -- CP-element group 52: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_408_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_Sample/rr
      -- 
    ca_1091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_408_inst_ack_1, ack => zeropad3D_CP_676_elements(52)); -- 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(52), ack => type_cast_412_inst_req_0); -- 
    rr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(52), ack => RPIPE_zeropad_input_pipe_426_inst_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_Sample/ra
      -- 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_412_inst_ack_0, ack => zeropad3D_CP_676_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	166 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	71 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_Update/ca
      -- 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_412_inst_ack_1, ack => zeropad3D_CP_676_elements(54)); -- 
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_update_start_
      -- CP-element group 55: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_Update/cr
      -- 
    ra_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_426_inst_ack_0, ack => zeropad3D_CP_676_elements(55)); -- 
    cr_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(55), ack => RPIPE_zeropad_input_pipe_426_inst_req_1); -- 
    -- CP-element group 56:  fork  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	59 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_426_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_Sample/rr
      -- 
    ca_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_426_inst_ack_1, ack => zeropad3D_CP_676_elements(56)); -- 
    rr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(56), ack => type_cast_430_inst_req_0); -- 
    rr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(56), ack => RPIPE_zeropad_input_pipe_444_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_Sample/ra
      -- 
    ra_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_430_inst_ack_0, ack => zeropad3D_CP_676_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	166 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	71 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_Update/ca
      -- 
    ca_1133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_430_inst_ack_1, ack => zeropad3D_CP_676_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	56 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_update_start_
      -- CP-element group 59: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_Sample/ra
      -- CP-element group 59: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_Update/cr
      -- 
    ra_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_444_inst_ack_0, ack => zeropad3D_CP_676_elements(59)); -- 
    cr_1146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(59), ack => RPIPE_zeropad_input_pipe_444_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	63 
    -- CP-element group 60:  members (9) 
      -- CP-element group 60: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_444_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_Sample/rr
      -- 
    ca_1147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_444_inst_ack_1, ack => zeropad3D_CP_676_elements(60)); -- 
    rr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(60), ack => type_cast_448_inst_req_0); -- 
    rr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(60), ack => RPIPE_zeropad_input_pipe_462_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_Sample/ra
      -- 
    ra_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_448_inst_ack_0, ack => zeropad3D_CP_676_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	166 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	71 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_Update/ca
      -- 
    ca_1161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_448_inst_ack_1, ack => zeropad3D_CP_676_elements(62)); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	60 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_update_start_
      -- CP-element group 63: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_Update/cr
      -- 
    ra_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_462_inst_ack_0, ack => zeropad3D_CP_676_elements(63)); -- 
    cr_1174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(63), ack => RPIPE_zeropad_input_pipe_462_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	67 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_462_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_Sample/rr
      -- 
    ca_1175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_462_inst_ack_1, ack => zeropad3D_CP_676_elements(64)); -- 
    rr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(64), ack => type_cast_466_inst_req_0); -- 
    rr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(64), ack => RPIPE_zeropad_input_pipe_480_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_Sample/ra
      -- 
    ra_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_466_inst_ack_0, ack => zeropad3D_CP_676_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	166 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	71 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_Update/ca
      -- 
    ca_1189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_466_inst_ack_1, ack => zeropad3D_CP_676_elements(66)); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	64 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_update_start_
      -- CP-element group 67: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_Update/cr
      -- 
    ra_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_480_inst_ack_0, ack => zeropad3D_CP_676_elements(67)); -- 
    cr_1202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(67), ack => RPIPE_zeropad_input_pipe_480_inst_req_1); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (6) 
      -- CP-element group 68: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_480_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_Sample/rr
      -- 
    ca_1203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_480_inst_ack_1, ack => zeropad3D_CP_676_elements(68)); -- 
    rr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(68), ack => type_cast_484_inst_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_Sample/ra
      -- 
    ra_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_484_inst_ack_0, ack => zeropad3D_CP_676_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	166 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_Update/ca
      -- 
    ca_1217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_484_inst_ack_1, ack => zeropad3D_CP_676_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	38 
    -- CP-element group 71: 	42 
    -- CP-element group 71: 	46 
    -- CP-element group 71: 	50 
    -- CP-element group 71: 	54 
    -- CP-element group 71: 	58 
    -- CP-element group 71: 	62 
    -- CP-element group 71: 	66 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/ptr_deref_492_Split/$entry
      -- CP-element group 71: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/ptr_deref_492_Split/$exit
      -- CP-element group 71: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/ptr_deref_492_Split/split_req
      -- CP-element group 71: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/ptr_deref_492_Split/split_ack
      -- CP-element group 71: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/word_access_start/$entry
      -- CP-element group 71: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/word_access_start/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/word_access_start/word_0/rr
      -- 
    rr_1255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(71), ack => ptr_deref_492_store_0_req_0); -- 
    zeropad3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(38) & zeropad3D_CP_676_elements(42) & zeropad3D_CP_676_elements(46) & zeropad3D_CP_676_elements(50) & zeropad3D_CP_676_elements(54) & zeropad3D_CP_676_elements(58) & zeropad3D_CP_676_elements(62) & zeropad3D_CP_676_elements(66) & zeropad3D_CP_676_elements(70);
      gj_zeropad3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/word_access_start/$exit
      -- CP-element group 72: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/word_access_start/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Sample/word_access_start/word_0/ra
      -- 
    ra_1256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_492_store_0_ack_0, ack => zeropad3D_CP_676_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	166 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Update/word_access_complete/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Update/word_access_complete/word_0/ca
      -- 
    ca_1267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_492_store_0_ack_1, ack => zeropad3D_CP_676_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	35 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_231/if_stmt_506__entry__
      -- CP-element group 74: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505__exit__
      -- CP-element group 74: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/$exit
      -- CP-element group 74: 	 branch_block_stmt_231/if_stmt_506_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_231/if_stmt_506_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_231/if_stmt_506_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_231/if_stmt_506_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_231/R_exitcond8_507_place
      -- CP-element group 74: 	 branch_block_stmt_231/if_stmt_506_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_231/if_stmt_506_else_link/$entry
      -- 
    branch_req_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(74), ack => if_stmt_506_branch_req_0); -- 
    zeropad3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(35) & zeropad3D_CP_676_elements(73);
      gj_zeropad3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  transition  place  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	167 
    -- CP-element group 75:  members (13) 
      -- CP-element group 75: 	 branch_block_stmt_231/forx_xendx_xloopexit_forx_xend
      -- CP-element group 75: 	 branch_block_stmt_231/merge_stmt_512__exit__
      -- CP-element group 75: 	 branch_block_stmt_231/if_stmt_506_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_231/if_stmt_506_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_231/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 75: 	 branch_block_stmt_231/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_231/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_231/merge_stmt_512_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_231/merge_stmt_512_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_231/merge_stmt_512_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_231/merge_stmt_512_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_231/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_231/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_506_branch_ack_1, ack => zeropad3D_CP_676_elements(75)); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	162 
    -- CP-element group 76: 	163 
    -- CP-element group 76:  members (12) 
      -- CP-element group 76: 	 branch_block_stmt_231/if_stmt_506_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_231/if_stmt_506_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_231/forx_xbody_forx_xbody
      -- CP-element group 76: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/$entry
      -- CP-element group 76: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/$entry
      -- CP-element group 76: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_506_branch_ack_0, ack => zeropad3D_CP_676_elements(76)); -- 
    rr_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(76), ack => type_cast_349_inst_req_0); -- 
    cr_1916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(76), ack => type_cast_349_inst_req_1); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	167 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_Sample/cra
      -- 
    cra_1298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_517_call_ack_0, ack => zeropad3D_CP_676_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	167 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_Update/cca
      -- CP-element group 78: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_Sample/rr
      -- 
    cca_1303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_517_call_ack_1, ack => zeropad3D_CP_676_elements(78)); -- 
    rr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(78), ack => type_cast_522_inst_req_0); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_Sample/ra
      -- 
    ra_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_522_inst_ack_0, ack => zeropad3D_CP_676_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	167 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	145 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_Update/ca
      -- 
    ca_1317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_522_inst_ack_1, ack => zeropad3D_CP_676_elements(80)); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	167 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_update_start_
      -- CP-element group 81: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_Sample/ack
      -- CP-element group 81: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_Update/req
      -- 
    ack_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_524_inst_ack_0, ack => zeropad3D_CP_676_elements(81)); -- 
    req_1330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(81), ack => WPIPE_Block0_starting_524_inst_req_1); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_Update/ack
      -- CP-element group 82: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_Sample/req
      -- 
    ack_1331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_524_inst_ack_1, ack => zeropad3D_CP_676_elements(82)); -- 
    req_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(82), ack => WPIPE_Block0_starting_527_inst_req_0); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_update_start_
      -- CP-element group 83: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_Sample/ack
      -- CP-element group 83: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_Update/req
      -- 
    ack_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_527_inst_ack_0, ack => zeropad3D_CP_676_elements(83)); -- 
    req_1344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(83), ack => WPIPE_Block0_starting_527_inst_req_1); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_527_Update/ack
      -- CP-element group 84: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_Sample/req
      -- 
    ack_1345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_527_inst_ack_1, ack => zeropad3D_CP_676_elements(84)); -- 
    req_1353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(84), ack => WPIPE_Block0_starting_530_inst_req_0); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_update_start_
      -- CP-element group 85: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_Sample/ack
      -- CP-element group 85: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_Update/req
      -- 
    ack_1354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_530_inst_ack_0, ack => zeropad3D_CP_676_elements(85)); -- 
    req_1358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(85), ack => WPIPE_Block0_starting_530_inst_req_1); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_530_Update/ack
      -- CP-element group 86: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_Sample/req
      -- 
    ack_1359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_530_inst_ack_1, ack => zeropad3D_CP_676_elements(86)); -- 
    req_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(86), ack => WPIPE_Block0_starting_533_inst_req_0); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_update_start_
      -- CP-element group 87: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_Update/req
      -- 
    ack_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_533_inst_ack_0, ack => zeropad3D_CP_676_elements(87)); -- 
    req_1372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(87), ack => WPIPE_Block0_starting_533_inst_req_1); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_533_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_Sample/req
      -- 
    ack_1373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_533_inst_ack_1, ack => zeropad3D_CP_676_elements(88)); -- 
    req_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(88), ack => WPIPE_Block0_starting_536_inst_req_0); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_update_start_
      -- CP-element group 89: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_Sample/ack
      -- CP-element group 89: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_Update/req
      -- 
    ack_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_536_inst_ack_0, ack => zeropad3D_CP_676_elements(89)); -- 
    req_1386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(89), ack => WPIPE_Block0_starting_536_inst_req_1); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_536_Update/ack
      -- CP-element group 90: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_Sample/req
      -- 
    ack_1387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_536_inst_ack_1, ack => zeropad3D_CP_676_elements(90)); -- 
    req_1395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(90), ack => WPIPE_Block0_starting_539_inst_req_0); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_update_start_
      -- CP-element group 91: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_Update/req
      -- 
    ack_1396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_539_inst_ack_0, ack => zeropad3D_CP_676_elements(91)); -- 
    req_1400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(91), ack => WPIPE_Block0_starting_539_inst_req_1); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_539_Update/ack
      -- CP-element group 92: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_Sample/req
      -- 
    ack_1401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_539_inst_ack_1, ack => zeropad3D_CP_676_elements(92)); -- 
    req_1409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(92), ack => WPIPE_Block0_starting_542_inst_req_0); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_update_start_
      -- CP-element group 93: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_Sample/ack
      -- CP-element group 93: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_Update/req
      -- 
    ack_1410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_542_inst_ack_0, ack => zeropad3D_CP_676_elements(93)); -- 
    req_1414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(93), ack => WPIPE_Block0_starting_542_inst_req_1); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	145 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_542_Update/ack
      -- 
    ack_1415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_542_inst_ack_1, ack => zeropad3D_CP_676_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	167 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_update_start_
      -- CP-element group 95: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_Sample/ack
      -- CP-element group 95: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_Update/req
      -- 
    ack_1424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_545_inst_ack_0, ack => zeropad3D_CP_676_elements(95)); -- 
    req_1428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(95), ack => WPIPE_Block1_starting_545_inst_req_1); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (6) 
      -- CP-element group 96: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_Update/ack
      -- CP-element group 96: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_Sample/req
      -- 
    ack_1429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_545_inst_ack_1, ack => zeropad3D_CP_676_elements(96)); -- 
    req_1437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(96), ack => WPIPE_Block1_starting_548_inst_req_0); -- 
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_Update/req
      -- CP-element group 97: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_update_start_
      -- CP-element group 97: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_Sample/ack
      -- 
    ack_1438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_548_inst_ack_0, ack => zeropad3D_CP_676_elements(97)); -- 
    req_1442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(97), ack => WPIPE_Block1_starting_548_inst_req_1); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_Sample/req
      -- CP-element group 98: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_Update/ack
      -- CP-element group 98: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_548_update_completed_
      -- 
    ack_1443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_548_inst_ack_1, ack => zeropad3D_CP_676_elements(98)); -- 
    req_1451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(98), ack => WPIPE_Block1_starting_551_inst_req_0); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_Sample/ack
      -- CP-element group 99: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_update_start_
      -- CP-element group 99: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_Update/req
      -- 
    ack_1452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_551_inst_ack_0, ack => zeropad3D_CP_676_elements(99)); -- 
    req_1456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(99), ack => WPIPE_Block1_starting_551_inst_req_1); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_Sample/req
      -- CP-element group 100: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_551_Update/ack
      -- 
    ack_1457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_551_inst_ack_1, ack => zeropad3D_CP_676_elements(100)); -- 
    req_1465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(100), ack => WPIPE_Block1_starting_554_inst_req_0); -- 
    -- CP-element group 101:  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_Update/req
      -- CP-element group 101: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_Sample/ack
      -- CP-element group 101: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_update_start_
      -- CP-element group 101: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_sample_completed_
      -- 
    ack_1466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_554_inst_ack_0, ack => zeropad3D_CP_676_elements(101)); -- 
    req_1470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(101), ack => WPIPE_Block1_starting_554_inst_req_1); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_Update/ack
      -- CP-element group 102: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_554_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_Sample/req
      -- 
    ack_1471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_554_inst_ack_1, ack => zeropad3D_CP_676_elements(102)); -- 
    req_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(102), ack => WPIPE_Block1_starting_557_inst_req_0); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_update_start_
      -- CP-element group 103: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_Update/req
      -- CP-element group 103: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_Sample/ack
      -- CP-element group 103: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_Sample/$exit
      -- 
    ack_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_557_inst_ack_0, ack => zeropad3D_CP_676_elements(103)); -- 
    req_1484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(103), ack => WPIPE_Block1_starting_557_inst_req_1); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (6) 
      -- CP-element group 104: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_Sample/req
      -- CP-element group 104: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_Update/ack
      -- CP-element group 104: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_557_Update/$exit
      -- 
    ack_1485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_557_inst_ack_1, ack => zeropad3D_CP_676_elements(104)); -- 
    req_1493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(104), ack => WPIPE_Block1_starting_560_inst_req_0); -- 
    -- CP-element group 105:  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (6) 
      -- CP-element group 105: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_Update/req
      -- CP-element group 105: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_Sample/ack
      -- CP-element group 105: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_update_start_
      -- CP-element group 105: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_sample_completed_
      -- 
    ack_1494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_560_inst_ack_0, ack => zeropad3D_CP_676_elements(105)); -- 
    req_1498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(105), ack => WPIPE_Block1_starting_560_inst_req_1); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_Sample/req
      -- CP-element group 106: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_Update/ack
      -- CP-element group 106: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_560_update_completed_
      -- 
    ack_1499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_560_inst_ack_1, ack => zeropad3D_CP_676_elements(106)); -- 
    req_1507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(106), ack => WPIPE_Block1_starting_563_inst_req_0); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_Update/req
      -- CP-element group 107: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_Sample/ack
      -- CP-element group 107: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_update_start_
      -- CP-element group 107: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_sample_completed_
      -- 
    ack_1508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_563_inst_ack_0, ack => zeropad3D_CP_676_elements(107)); -- 
    req_1512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(107), ack => WPIPE_Block1_starting_563_inst_req_1); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	145 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_Update/ack
      -- CP-element group 108: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_563_update_completed_
      -- 
    ack_1513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_starting_563_inst_ack_1, ack => zeropad3D_CP_676_elements(108)); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	167 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_Sample/ack
      -- CP-element group 109: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_update_start_
      -- CP-element group 109: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_Update/req
      -- CP-element group 109: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_Sample/$exit
      -- 
    ack_1522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_566_inst_ack_0, ack => zeropad3D_CP_676_elements(109)); -- 
    req_1526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(109), ack => WPIPE_Block2_starting_566_inst_req_1); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_Update/ack
      -- CP-element group 110: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_Sample/req
      -- CP-element group 110: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_sample_start_
      -- 
    ack_1527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_566_inst_ack_1, ack => zeropad3D_CP_676_elements(110)); -- 
    req_1535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(110), ack => WPIPE_Block2_starting_569_inst_req_0); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_Update/req
      -- CP-element group 111: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_Sample/ack
      -- CP-element group 111: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_update_start_
      -- CP-element group 111: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_sample_completed_
      -- 
    ack_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_569_inst_ack_0, ack => zeropad3D_CP_676_elements(111)); -- 
    req_1540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => WPIPE_Block2_starting_569_inst_req_1); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (6) 
      -- CP-element group 112: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_Update/ack
      -- CP-element group 112: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_Sample/req
      -- CP-element group 112: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_569_update_completed_
      -- 
    ack_1541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_569_inst_ack_1, ack => zeropad3D_CP_676_elements(112)); -- 
    req_1549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(112), ack => WPIPE_Block2_starting_572_inst_req_0); -- 
    -- CP-element group 113:  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (6) 
      -- CP-element group 113: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_Sample/ack
      -- CP-element group 113: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_update_start_
      -- CP-element group 113: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_Update/req
      -- 
    ack_1550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_572_inst_ack_0, ack => zeropad3D_CP_676_elements(113)); -- 
    req_1554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(113), ack => WPIPE_Block2_starting_572_inst_req_1); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_Sample/req
      -- CP-element group 114: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_Update/ack
      -- CP-element group 114: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_572_Update/$exit
      -- 
    ack_1555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_572_inst_ack_1, ack => zeropad3D_CP_676_elements(114)); -- 
    req_1563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(114), ack => WPIPE_Block2_starting_575_inst_req_0); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_Update/req
      -- CP-element group 115: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_Sample/ack
      -- CP-element group 115: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_update_start_
      -- CP-element group 115: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_sample_completed_
      -- 
    ack_1564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_575_inst_ack_0, ack => zeropad3D_CP_676_elements(115)); -- 
    req_1568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(115), ack => WPIPE_Block2_starting_575_inst_req_1); -- 
    -- CP-element group 116:  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (6) 
      -- CP-element group 116: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_Sample/req
      -- CP-element group 116: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_Update/ack
      -- CP-element group 116: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_575_update_completed_
      -- 
    ack_1569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_575_inst_ack_1, ack => zeropad3D_CP_676_elements(116)); -- 
    req_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(116), ack => WPIPE_Block2_starting_578_inst_req_0); -- 
    -- CP-element group 117:  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (6) 
      -- CP-element group 117: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_Update/req
      -- CP-element group 117: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_Sample/ack
      -- CP-element group 117: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_update_start_
      -- CP-element group 117: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_sample_completed_
      -- 
    ack_1578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_578_inst_ack_0, ack => zeropad3D_CP_676_elements(117)); -- 
    req_1582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(117), ack => WPIPE_Block2_starting_578_inst_req_1); -- 
    -- CP-element group 118:  transition  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (6) 
      -- CP-element group 118: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_Sample/req
      -- CP-element group 118: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_Update/ack
      -- CP-element group 118: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_578_update_completed_
      -- 
    ack_1583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_578_inst_ack_1, ack => zeropad3D_CP_676_elements(118)); -- 
    req_1591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(118), ack => WPIPE_Block2_starting_581_inst_req_0); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_Update/req
      -- CP-element group 119: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_Sample/ack
      -- CP-element group 119: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_update_start_
      -- CP-element group 119: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_sample_completed_
      -- 
    ack_1592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_581_inst_ack_0, ack => zeropad3D_CP_676_elements(119)); -- 
    req_1596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(119), ack => WPIPE_Block2_starting_581_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_Sample/req
      -- CP-element group 120: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_Update/ack
      -- CP-element group 120: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_581_update_completed_
      -- 
    ack_1597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_581_inst_ack_1, ack => zeropad3D_CP_676_elements(120)); -- 
    req_1605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(120), ack => WPIPE_Block2_starting_584_inst_req_0); -- 
    -- CP-element group 121:  transition  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (6) 
      -- CP-element group 121: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_Sample/ack
      -- CP-element group 121: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_update_start_
      -- CP-element group 121: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_Update/req
      -- CP-element group 121: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_sample_completed_
      -- 
    ack_1606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_584_inst_ack_0, ack => zeropad3D_CP_676_elements(121)); -- 
    req_1610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(121), ack => WPIPE_Block2_starting_584_inst_req_1); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	145 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_Update/ack
      -- CP-element group 122: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_584_Update/$exit
      -- 
    ack_1611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_starting_584_inst_ack_1, ack => zeropad3D_CP_676_elements(122)); -- 
    -- CP-element group 123:  transition  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	167 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (6) 
      -- CP-element group 123: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_Sample/ack
      -- CP-element group 123: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_update_start_
      -- CP-element group 123: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_Update/req
      -- 
    ack_1620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_587_inst_ack_0, ack => zeropad3D_CP_676_elements(123)); -- 
    req_1624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(123), ack => WPIPE_Block3_starting_587_inst_req_1); -- 
    -- CP-element group 124:  transition  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (6) 
      -- CP-element group 124: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_Update/ack
      -- CP-element group 124: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_Sample/req
      -- CP-element group 124: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_sample_start_
      -- 
    ack_1625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_587_inst_ack_1, ack => zeropad3D_CP_676_elements(124)); -- 
    req_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => WPIPE_Block3_starting_590_inst_req_0); -- 
    -- CP-element group 125:  transition  input  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (6) 
      -- CP-element group 125: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_Update/req
      -- CP-element group 125: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_Update/$entry
      -- CP-element group 125: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_Sample/ack
      -- CP-element group 125: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_update_start_
      -- CP-element group 125: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_sample_completed_
      -- 
    ack_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_590_inst_ack_0, ack => zeropad3D_CP_676_elements(125)); -- 
    req_1638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(125), ack => WPIPE_Block3_starting_590_inst_req_1); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (6) 
      -- CP-element group 126: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_Sample/req
      -- CP-element group 126: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_590_update_completed_
      -- 
    ack_1639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_590_inst_ack_1, ack => zeropad3D_CP_676_elements(126)); -- 
    req_1647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(126), ack => WPIPE_Block3_starting_593_inst_req_0); -- 
    -- CP-element group 127:  transition  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (6) 
      -- CP-element group 127: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_Update/req
      -- CP-element group 127: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_Sample/ack
      -- CP-element group 127: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_update_start_
      -- CP-element group 127: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_Update/$entry
      -- 
    ack_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_593_inst_ack_0, ack => zeropad3D_CP_676_elements(127)); -- 
    req_1652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(127), ack => WPIPE_Block3_starting_593_inst_req_1); -- 
    -- CP-element group 128:  transition  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (6) 
      -- CP-element group 128: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_Update/ack
      -- CP-element group 128: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_Sample/req
      -- CP-element group 128: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_593_Update/$exit
      -- 
    ack_1653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_593_inst_ack_1, ack => zeropad3D_CP_676_elements(128)); -- 
    req_1661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => WPIPE_Block3_starting_596_inst_req_0); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_update_start_
      -- CP-element group 129: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_Sample/ack
      -- CP-element group 129: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_Update/req
      -- CP-element group 129: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_Update/$entry
      -- 
    ack_1662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_596_inst_ack_0, ack => zeropad3D_CP_676_elements(129)); -- 
    req_1666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(129), ack => WPIPE_Block3_starting_596_inst_req_1); -- 
    -- CP-element group 130:  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (6) 
      -- CP-element group 130: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_Sample/req
      -- CP-element group 130: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_Update/ack
      -- CP-element group 130: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_596_Update/$exit
      -- 
    ack_1667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_596_inst_ack_1, ack => zeropad3D_CP_676_elements(130)); -- 
    req_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(130), ack => WPIPE_Block3_starting_599_inst_req_0); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_Update/req
      -- CP-element group 131: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_Sample/ack
      -- CP-element group 131: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_update_start_
      -- CP-element group 131: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_sample_completed_
      -- 
    ack_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_599_inst_ack_0, ack => zeropad3D_CP_676_elements(131)); -- 
    req_1680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(131), ack => WPIPE_Block3_starting_599_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_Sample/req
      -- CP-element group 132: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_Update/ack
      -- CP-element group 132: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_599_update_completed_
      -- 
    ack_1681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_599_inst_ack_1, ack => zeropad3D_CP_676_elements(132)); -- 
    req_1689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(132), ack => WPIPE_Block3_starting_602_inst_req_0); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_Update/req
      -- CP-element group 133: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_Sample/ack
      -- CP-element group 133: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_update_start_
      -- 
    ack_1690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_602_inst_ack_0, ack => zeropad3D_CP_676_elements(133)); -- 
    req_1694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(133), ack => WPIPE_Block3_starting_602_inst_req_1); -- 
    -- CP-element group 134:  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_Update/ack
      -- CP-element group 134: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_602_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_Sample/req
      -- CP-element group 134: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_Sample/$entry
      -- 
    ack_1695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_602_inst_ack_1, ack => zeropad3D_CP_676_elements(134)); -- 
    req_1703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(134), ack => WPIPE_Block3_starting_605_inst_req_0); -- 
    -- CP-element group 135:  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (6) 
      -- CP-element group 135: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_Update/req
      -- CP-element group 135: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_Sample/ack
      -- CP-element group 135: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_update_start_
      -- CP-element group 135: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_sample_completed_
      -- 
    ack_1704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_605_inst_ack_0, ack => zeropad3D_CP_676_elements(135)); -- 
    req_1708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(135), ack => WPIPE_Block3_starting_605_inst_req_1); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	145 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_Update/ack
      -- CP-element group 136: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_605_update_completed_
      -- 
    ack_1709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_starting_605_inst_ack_1, ack => zeropad3D_CP_676_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	167 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_Update/cr
      -- CP-element group 137: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_update_start_
      -- CP-element group 137: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_sample_completed_
      -- 
    ra_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_complete_609_inst_ack_0, ack => zeropad3D_CP_676_elements(137)); -- 
    cr_1722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(137), ack => RPIPE_Block0_complete_609_inst_req_1); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	145 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_update_completed_
      -- 
    ca_1723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_complete_609_inst_ack_1, ack => zeropad3D_CP_676_elements(138)); -- 
    -- CP-element group 139:  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	167 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139:  members (6) 
      -- CP-element group 139: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_Update/cr
      -- CP-element group 139: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_Sample/ra
      -- CP-element group 139: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_update_start_
      -- CP-element group 139: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_sample_completed_
      -- 
    ra_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_complete_612_inst_ack_0, ack => zeropad3D_CP_676_elements(139)); -- 
    cr_1736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(139), ack => RPIPE_Block1_complete_612_inst_req_1); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	145 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_update_completed_
      -- 
    ca_1737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_complete_612_inst_ack_1, ack => zeropad3D_CP_676_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	167 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_update_start_
      -- CP-element group 141: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_Update/cr
      -- 
    ra_1746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_complete_615_inst_ack_0, ack => zeropad3D_CP_676_elements(141)); -- 
    cr_1750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(141), ack => RPIPE_Block2_complete_615_inst_req_1); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_Update/$exit
      -- 
    ca_1751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_complete_615_inst_ack_1, ack => zeropad3D_CP_676_elements(142)); -- 
    -- CP-element group 143:  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	167 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (6) 
      -- CP-element group 143: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_update_start_
      -- CP-element group 143: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_Update/cr
      -- CP-element group 143: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_Sample/$exit
      -- 
    ra_1760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_complete_618_inst_ack_0, ack => zeropad3D_CP_676_elements(143)); -- 
    cr_1764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(143), ack => RPIPE_Block3_complete_618_inst_req_1); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_Update/$exit
      -- 
    ca_1765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_complete_618_inst_ack_1, ack => zeropad3D_CP_676_elements(144)); -- 
    -- CP-element group 145:  join  fork  transition  place  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	80 
    -- CP-element group 145: 	94 
    -- CP-element group 145: 	108 
    -- CP-element group 145: 	122 
    -- CP-element group 145: 	136 
    -- CP-element group 145: 	138 
    -- CP-element group 145: 	140 
    -- CP-element group 145: 	142 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145: 	147 
    -- CP-element group 145: 	149 
    -- CP-element group 145:  members (13) 
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619__exit__
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635__entry__
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_update_start_
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_Update/ccr
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_Sample/crr
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_update_start_
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/$entry
      -- CP-element group 145: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/$exit
      -- 
    cr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(145), ack => type_cast_626_inst_req_1); -- 
    ccr_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(145), ack => call_stmt_622_call_req_1); -- 
    crr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(145), ack => call_stmt_622_call_req_0); -- 
    zeropad3D_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(80) & zeropad3D_CP_676_elements(94) & zeropad3D_CP_676_elements(108) & zeropad3D_CP_676_elements(122) & zeropad3D_CP_676_elements(136) & zeropad3D_CP_676_elements(138) & zeropad3D_CP_676_elements(140) & zeropad3D_CP_676_elements(142) & zeropad3D_CP_676_elements(144);
      gj_zeropad3D_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_Sample/cra
      -- CP-element group 146: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_sample_completed_
      -- 
    cra_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_622_call_ack_0, ack => zeropad3D_CP_676_elements(146)); -- 
    -- CP-element group 147:  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (6) 
      -- CP-element group 147: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_Update/cca
      -- CP-element group 147: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/call_stmt_622_update_completed_
      -- 
    cca_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_622_call_ack_1, ack => zeropad3D_CP_676_elements(147)); -- 
    rr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(147), ack => type_cast_626_inst_req_0); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_Sample/ra
      -- 
    ra_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_626_inst_ack_0, ack => zeropad3D_CP_676_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	145 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/type_cast_626_Update/ca
      -- CP-element group 149: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_Sample/req
      -- CP-element group 149: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_sample_start_
      -- 
    ca_1796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_626_inst_ack_1, ack => zeropad3D_CP_676_elements(149)); -- 
    req_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(149), ack => WPIPE_elapsed_time_pipe_633_inst_req_0); -- 
    -- CP-element group 150:  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (6) 
      -- CP-element group 150: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_Update/req
      -- CP-element group 150: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_Sample/ack
      -- CP-element group 150: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_update_start_
      -- CP-element group 150: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_sample_completed_
      -- 
    ack_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_633_inst_ack_0, ack => zeropad3D_CP_676_elements(150)); -- 
    req_1809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(150), ack => WPIPE_elapsed_time_pipe_633_inst_req_1); -- 
    -- CP-element group 151:  fork  transition  place  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: 	153 
    -- CP-element group 151: 	154 
    -- CP-element group 151: 	155 
    -- CP-element group 151: 	156 
    -- CP-element group 151: 	157 
    -- CP-element group 151: 	160 
    -- CP-element group 151:  members (28) 
      -- CP-element group 151: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_Update/ack
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_Update/cr
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660__entry__
      -- CP-element group 151: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635__exit__
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_Update/ccr
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/$entry
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_Update/cr
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_update_start_
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_update_start_
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/WPIPE_elapsed_time_pipe_633_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_231/call_stmt_622_to_assign_stmt_635/$exit
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_update_start_
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_Update/cr
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_update_start_
      -- 
    ack_1810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_633_inst_ack_1, ack => zeropad3D_CP_676_elements(151)); -- 
    cr_1840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(151), ack => type_cast_643_inst_req_1); -- 
    rr_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(151), ack => type_cast_643_inst_req_0); -- 
    ccr_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(151), ack => call_stmt_660_call_req_1); -- 
    cr_1854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(151), ack => type_cast_647_inst_req_1); -- 
    rr_1849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(151), ack => type_cast_647_inst_req_0); -- 
    cr_1826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(151), ack => type_cast_639_inst_req_1); -- 
    rr_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(151), ack => type_cast_639_inst_req_0); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_Sample/$exit
      -- 
    ra_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_639_inst_ack_0, ack => zeropad3D_CP_676_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	158 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_639_update_completed_
      -- 
    ca_1827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_639_inst_ack_1, ack => zeropad3D_CP_676_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	151 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_sample_completed_
      -- 
    ra_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_0, ack => zeropad3D_CP_676_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	151 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	158 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_643_Update/ca
      -- 
    ca_1841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_1, ack => zeropad3D_CP_676_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	151 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_sample_completed_
      -- 
    ra_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_647_inst_ack_0, ack => zeropad3D_CP_676_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	151 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/type_cast_647_update_completed_
      -- 
    ca_1855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_647_inst_ack_1, ack => zeropad3D_CP_676_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	153 
    -- CP-element group 158: 	155 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_Sample/crr
      -- 
    crr_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(158), ack => call_stmt_660_call_req_0); -- 
    zeropad3D_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(153) & zeropad3D_CP_676_elements(155) & zeropad3D_CP_676_elements(157);
      gj_zeropad3D_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_Sample/cra
      -- CP-element group 159: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_Sample/$exit
      -- 
    cra_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_660_call_ack_0, ack => zeropad3D_CP_676_elements(159)); -- 
    -- CP-element group 160:  transition  place  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	151 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (16) 
      -- CP-element group 160: 	 $exit
      -- CP-element group 160: 	 branch_block_stmt_231/branch_block_stmt_231__exit__
      -- CP-element group 160: 	 branch_block_stmt_231/merge_stmt_662__exit__
      -- CP-element group 160: 	 branch_block_stmt_231/return__
      -- CP-element group 160: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660__exit__
      -- CP-element group 160: 	 branch_block_stmt_231/$exit
      -- CP-element group 160: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/$exit
      -- CP-element group 160: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_231/assign_stmt_640_to_call_stmt_660/call_stmt_660_Update/cca
      -- CP-element group 160: 	 branch_block_stmt_231/return___PhiReq/$entry
      -- CP-element group 160: 	 branch_block_stmt_231/return___PhiReq/$exit
      -- CP-element group 160: 	 branch_block_stmt_231/merge_stmt_662_PhiReqMerge
      -- CP-element group 160: 	 branch_block_stmt_231/merge_stmt_662_PhiAck/$entry
      -- CP-element group 160: 	 branch_block_stmt_231/merge_stmt_662_PhiAck/$exit
      -- CP-element group 160: 	 branch_block_stmt_231/merge_stmt_662_PhiAck/dummy
      -- 
    cca_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_660_call_ack_1, ack => zeropad3D_CP_676_elements(160)); -- 
    -- CP-element group 161:  transition  output  delay-element  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	34 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	165 
    -- CP-element group 161:  members (5) 
      -- CP-element group 161: 	 branch_block_stmt_231/bbx_xnph_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_347_konst_delay_trans
      -- CP-element group 161: 	 branch_block_stmt_231/bbx_xnph_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/$exit
      -- CP-element group 161: 	 branch_block_stmt_231/bbx_xnph_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_req
      -- CP-element group 161: 	 branch_block_stmt_231/bbx_xnph_forx_xbody_PhiReq/phi_stmt_343/$exit
      -- CP-element group 161: 	 branch_block_stmt_231/bbx_xnph_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_343_req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_343_req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(161), ack => phi_stmt_343_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(161) is a control-delay.
    cp_element_161_delay: control_delay_element  generic map(name => " 161_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(34), ack => zeropad3D_CP_676_elements(161), clk => clk, reset =>reset);
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	76 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/SplitProtocol/Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/SplitProtocol/Sample/ra
      -- 
    ra_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_349_inst_ack_0, ack => zeropad3D_CP_676_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	76 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/SplitProtocol/Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/SplitProtocol/Update/ca
      -- 
    ca_1917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_349_inst_ack_1, ack => zeropad3D_CP_676_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (6) 
      -- CP-element group 164: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 164: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/$exit
      -- CP-element group 164: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/$exit
      -- CP-element group 164: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/$exit
      -- CP-element group 164: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_sources/type_cast_349/SplitProtocol/$exit
      -- CP-element group 164: 	 branch_block_stmt_231/forx_xbody_forx_xbody_PhiReq/phi_stmt_343/phi_stmt_343_req
      -- 
    phi_stmt_343_req_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_343_req_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(164), ack => phi_stmt_343_req_1); -- 
    zeropad3D_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(162) & zeropad3D_CP_676_elements(163);
      gj_zeropad3D_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	161 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_231/merge_stmt_342_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_231/merge_stmt_342_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(165) <= OrReduce(zeropad3D_CP_676_elements(161) & zeropad3D_CP_676_elements(164));
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	35 
    -- CP-element group 166: 	36 
    -- CP-element group 166: 	38 
    -- CP-element group 166: 	39 
    -- CP-element group 166: 	42 
    -- CP-element group 166: 	46 
    -- CP-element group 166: 	50 
    -- CP-element group 166: 	54 
    -- CP-element group 166: 	58 
    -- CP-element group 166: 	62 
    -- CP-element group 166: 	66 
    -- CP-element group 166: 	70 
    -- CP-element group 166: 	73 
    -- CP-element group 166:  members (56) 
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505__entry__
      -- CP-element group 166: 	 branch_block_stmt_231/merge_stmt_342__exit__
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_update_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_resized_1
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_scaled_1
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_computed_1
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_resize_1/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_resize_1/$exit
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_resize_1/index_resize_req
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_resize_1/index_resize_ack
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_scale_1/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_scale_1/$exit
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_scale_1/scale_rename_req
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_index_scale_1/scale_rename_ack
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_final_index_sum_regn_update_start
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_final_index_sum_regn_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_final_index_sum_regn_Sample/req
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_final_index_sum_regn_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/array_obj_ref_355_final_index_sum_regn_Update/req
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_complete/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/addr_of_356_complete/req
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/RPIPE_zeropad_input_pipe_359_Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_update_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_363_Update/cr
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_update_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_376_Update/cr
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_update_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_394_Update/cr
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_update_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_412_Update/cr
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_update_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_430_Update/cr
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_update_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_448_Update/cr
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_update_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_466_Update/cr
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_update_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/type_cast_484_Update/cr
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_update_start_
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Update/word_access_complete/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Update/word_access_complete/word_0/$entry
      -- CP-element group 166: 	 branch_block_stmt_231/assign_stmt_357_to_assign_stmt_505/ptr_deref_492_Update/word_access_complete/word_0/cr
      -- CP-element group 166: 	 branch_block_stmt_231/merge_stmt_342_PhiAck/$exit
      -- CP-element group 166: 	 branch_block_stmt_231/merge_stmt_342_PhiAck/phi_stmt_343_ack
      -- 
    phi_stmt_343_ack_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_343_ack_0, ack => zeropad3D_CP_676_elements(166)); -- 
    req_972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => array_obj_ref_355_index_offset_req_0); -- 
    req_977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => array_obj_ref_355_index_offset_req_1); -- 
    req_992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => addr_of_356_final_reg_req_1); -- 
    rr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => RPIPE_zeropad_input_pipe_359_inst_req_0); -- 
    cr_1020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => type_cast_363_inst_req_1); -- 
    cr_1048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => type_cast_376_inst_req_1); -- 
    cr_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => type_cast_394_inst_req_1); -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => type_cast_412_inst_req_1); -- 
    cr_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => type_cast_430_inst_req_1); -- 
    cr_1160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => type_cast_448_inst_req_1); -- 
    cr_1188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => type_cast_466_inst_req_1); -- 
    cr_1216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => type_cast_484_inst_req_1); -- 
    cr_1266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => ptr_deref_492_store_0_req_1); -- 
    -- CP-element group 167:  merge  fork  transition  place  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	26 
    -- CP-element group 167: 	75 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	77 
    -- CP-element group 167: 	78 
    -- CP-element group 167: 	80 
    -- CP-element group 167: 	81 
    -- CP-element group 167: 	95 
    -- CP-element group 167: 	109 
    -- CP-element group 167: 	123 
    -- CP-element group 167: 	137 
    -- CP-element group 167: 	139 
    -- CP-element group 167: 	141 
    -- CP-element group 167: 	143 
    -- CP-element group 167:  members (40) 
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_Sample/req
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_Sample/req
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619__entry__
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/merge_stmt_514__exit__
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block2_starting_566_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block3_starting_587_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block2_complete_615_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block0_complete_609_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block1_complete_612_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_update_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_Sample/crr
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/call_stmt_517_Update/ccr
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_update_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/RPIPE_Block3_complete_618_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/type_cast_522_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block0_starting_524_Sample/req
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/call_stmt_517_to_assign_stmt_619/WPIPE_Block1_starting_545_Sample/req
      -- CP-element group 167: 	 branch_block_stmt_231/merge_stmt_514_PhiReqMerge
      -- CP-element group 167: 	 branch_block_stmt_231/merge_stmt_514_PhiAck/$entry
      -- CP-element group 167: 	 branch_block_stmt_231/merge_stmt_514_PhiAck/$exit
      -- CP-element group 167: 	 branch_block_stmt_231/merge_stmt_514_PhiAck/dummy
      -- 
    req_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => WPIPE_Block2_starting_566_inst_req_0); -- 
    req_1619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => WPIPE_Block3_starting_587_inst_req_0); -- 
    rr_1717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => RPIPE_Block0_complete_609_inst_req_0); -- 
    rr_1745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => RPIPE_Block2_complete_615_inst_req_0); -- 
    rr_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => RPIPE_Block1_complete_612_inst_req_0); -- 
    crr_1297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => call_stmt_517_call_req_0); -- 
    rr_1759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => RPIPE_Block3_complete_618_inst_req_0); -- 
    ccr_1302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => call_stmt_517_call_req_1); -- 
    cr_1316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => type_cast_522_inst_req_1); -- 
    req_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => WPIPE_Block0_starting_524_inst_req_0); -- 
    req_1423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => WPIPE_Block1_starting_545_inst_req_0); -- 
    zeropad3D_CP_676_elements(167) <= OrReduce(zeropad3D_CP_676_elements(26) & zeropad3D_CP_676_elements(75));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_354_resized : std_logic_vector(13 downto 0);
    signal R_indvar_354_scaled : std_logic_vector(13 downto 0);
    signal add31_400 : std_logic_vector(63 downto 0);
    signal add37_418 : std_logic_vector(63 downto 0);
    signal add43_436 : std_logic_vector(63 downto 0);
    signal add49_454 : std_logic_vector(63 downto 0);
    signal add55_472 : std_logic_vector(63 downto 0);
    signal add61_490 : std_logic_vector(63 downto 0);
    signal add_382 : std_logic_vector(63 downto 0);
    signal array_obj_ref_355_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_355_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_355_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_355_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_355_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_355_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_357 : std_logic_vector(31 downto 0);
    signal call100_613 : std_logic_vector(7 downto 0);
    signal call103_616 : std_logic_vector(7 downto 0);
    signal call106_619 : std_logic_vector(7 downto 0);
    signal call109_622 : std_logic_vector(63 downto 0);
    signal call1_237 : std_logic_vector(7 downto 0);
    signal call20_360 : std_logic_vector(7 downto 0);
    signal call23_373 : std_logic_vector(7 downto 0);
    signal call28_391 : std_logic_vector(7 downto 0);
    signal call2_240 : std_logic_vector(7 downto 0);
    signal call34_409 : std_logic_vector(7 downto 0);
    signal call3_243 : std_logic_vector(7 downto 0);
    signal call40_427 : std_logic_vector(7 downto 0);
    signal call46_445 : std_logic_vector(7 downto 0);
    signal call4_246 : std_logic_vector(7 downto 0);
    signal call52_463 : std_logic_vector(7 downto 0);
    signal call58_481 : std_logic_vector(7 downto 0);
    signal call5_249 : std_logic_vector(7 downto 0);
    signal call66_517 : std_logic_vector(63 downto 0);
    signal call6_252 : std_logic_vector(7 downto 0);
    signal call7_255 : std_logic_vector(7 downto 0);
    signal call8_258 : std_logic_vector(7 downto 0);
    signal call97_610 : std_logic_vector(7 downto 0);
    signal call_234 : std_logic_vector(7 downto 0);
    signal cmp126_292 : std_logic_vector(0 downto 0);
    signal conv10_266 : std_logic_vector(63 downto 0);
    signal conv110_627 : std_logic_vector(63 downto 0);
    signal conv116_640 : std_logic_vector(31 downto 0);
    signal conv118_644 : std_logic_vector(31 downto 0);
    signal conv121_648 : std_logic_vector(31 downto 0);
    signal conv12_270 : std_logic_vector(63 downto 0);
    signal conv21_364 : std_logic_vector(63 downto 0);
    signal conv25_377 : std_logic_vector(63 downto 0);
    signal conv30_395 : std_logic_vector(63 downto 0);
    signal conv36_413 : std_logic_vector(63 downto 0);
    signal conv42_431 : std_logic_vector(63 downto 0);
    signal conv48_449 : std_logic_vector(63 downto 0);
    signal conv54_467 : std_logic_vector(63 downto 0);
    signal conv60_485 : std_logic_vector(63 downto 0);
    signal conv67_523 : std_logic_vector(63 downto 0);
    signal conv_262 : std_logic_vector(63 downto 0);
    signal exitcond8_505 : std_logic_vector(0 downto 0);
    signal indvar_343 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_500 : std_logic_vector(63 downto 0);
    signal mul119_653 : std_logic_vector(31 downto 0);
    signal mul122_658 : std_logic_vector(31 downto 0);
    signal mul13_280 : std_logic_vector(63 downto 0);
    signal mul_275 : std_logic_vector(63 downto 0);
    signal ptr_deref_492_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_492_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_492_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_492_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_492_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_492_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl27_388 : std_logic_vector(63 downto 0);
    signal shl33_406 : std_logic_vector(63 downto 0);
    signal shl39_424 : std_logic_vector(63 downto 0);
    signal shl45_442 : std_logic_vector(63 downto 0);
    signal shl51_460 : std_logic_vector(63 downto 0);
    signal shl57_478 : std_logic_vector(63 downto 0);
    signal shl_370 : std_logic_vector(63 downto 0);
    signal shr125x_xmask_286 : std_logic_vector(63 downto 0);
    signal sub_632 : std_logic_vector(63 downto 0);
    signal tmp1_307 : std_logic_vector(63 downto 0);
    signal tmp2_312 : std_logic_vector(63 downto 0);
    signal tmp3_316 : std_logic_vector(63 downto 0);
    signal tmp4_321 : std_logic_vector(63 downto 0);
    signal tmp5_327 : std_logic_vector(63 downto 0);
    signal tmp6_333 : std_logic_vector(0 downto 0);
    signal tmp_303 : std_logic_vector(63 downto 0);
    signal type_cast_284_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_290_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_325_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_331_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_338_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_347_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_349_wire : std_logic_vector(63 downto 0);
    signal type_cast_368_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_386_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_404_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_422_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_440_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_458_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_476_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_498_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_521_wire : std_logic_vector(63 downto 0);
    signal type_cast_625_wire : std_logic_vector(63 downto 0);
    signal umax7_340 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_355_constant_part_of_offset <= "00000000000000";
    array_obj_ref_355_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_355_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_355_resized_base_address <= "00000000000000";
    ptr_deref_492_word_offset_0 <= "00000000000000";
    type_cast_284_wire_constant <= "0000000000000000000000000000000000000000111111111111111111111100";
    type_cast_290_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_325_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_331_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_338_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_347_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_368_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_404_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_422_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_440_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_458_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_476_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_498_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_343: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_347_wire_constant & type_cast_349_wire;
      req <= phi_stmt_343_req_0 & phi_stmt_343_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_343",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_343_ack_0,
          idata => idata,
          odata => indvar_343,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_343
    -- flow-through select operator MUX_339_inst
    umax7_340 <= tmp5_327 when (tmp6_333(0) /=  '0') else type_cast_338_wire_constant;
    addr_of_356_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_356_final_reg_req_0;
      addr_of_356_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_356_final_reg_req_1;
      addr_of_356_final_reg_ack_1<= rack(0);
      addr_of_356_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_356_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_355_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_357,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_261_inst_req_0;
      type_cast_261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_261_inst_req_1;
      type_cast_261_inst_ack_1<= rack(0);
      type_cast_261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_265_inst_req_0;
      type_cast_265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_265_inst_req_1;
      type_cast_265_inst_ack_1<= rack(0);
      type_cast_265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_243,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_269_inst_req_0;
      type_cast_269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_269_inst_req_1;
      type_cast_269_inst_ack_1<= rack(0);
      type_cast_269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_302_inst_req_0;
      type_cast_302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_302_inst_req_1;
      type_cast_302_inst_ack_1<= rack(0);
      type_cast_302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_243,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp_303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_306_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_306_inst_req_0;
      type_cast_306_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_306_inst_req_1;
      type_cast_306_inst_ack_1<= rack(0);
      type_cast_306_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_306_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_307,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_315_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_315_inst_req_0;
      type_cast_315_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_315_inst_req_1;
      type_cast_315_inst_ack_1<= rack(0);
      type_cast_315_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_315_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_316,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_349_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_349_inst_req_0;
      type_cast_349_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_349_inst_req_1;
      type_cast_349_inst_ack_1<= rack(0);
      type_cast_349_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_349_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_349_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_363_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_363_inst_req_0;
      type_cast_363_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_363_inst_req_1;
      type_cast_363_inst_ack_1<= rack(0);
      type_cast_363_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_363_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_360,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv21_364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_376_inst_req_0;
      type_cast_376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_376_inst_req_1;
      type_cast_376_inst_ack_1<= rack(0);
      type_cast_376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_376_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv25_377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_394_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_394_inst_req_0;
      type_cast_394_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_394_inst_req_1;
      type_cast_394_inst_ack_1<= rack(0);
      type_cast_394_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_394_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_395,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_412_inst_req_0;
      type_cast_412_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_412_inst_req_1;
      type_cast_412_inst_ack_1<= rack(0);
      type_cast_412_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_412_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call34_409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_430_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_430_inst_req_0;
      type_cast_430_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_430_inst_req_1;
      type_cast_430_inst_ack_1<= rack(0);
      type_cast_430_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_430_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call40_427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_431,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_448_inst_req_0;
      type_cast_448_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_448_inst_req_1;
      type_cast_448_inst_ack_1<= rack(0);
      type_cast_448_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_448_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_445,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_449,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_466_inst_req_0;
      type_cast_466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_466_inst_req_1;
      type_cast_466_inst_ack_1<= rack(0);
      type_cast_466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call52_463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv54_467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_484_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_484_inst_req_0;
      type_cast_484_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_484_inst_req_1;
      type_cast_484_inst_ack_1<= rack(0);
      type_cast_484_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_484_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call58_481,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_485,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_522_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_522_inst_req_0;
      type_cast_522_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_522_inst_req_1;
      type_cast_522_inst_ack_1<= rack(0);
      type_cast_522_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_522_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_521_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_523,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_626_inst_req_0;
      type_cast_626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_626_inst_req_1;
      type_cast_626_inst_ack_1<= rack(0);
      type_cast_626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_625_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_627,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_639_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_639_inst_req_0;
      type_cast_639_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_639_inst_req_1;
      type_cast_639_inst_ack_1<= rack(0);
      type_cast_639_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_639_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_640,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_643_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_643_inst_req_0;
      type_cast_643_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_643_inst_req_1;
      type_cast_643_inst_ack_1<= rack(0);
      type_cast_643_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_643_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv118_644,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_647_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_647_inst_req_0;
      type_cast_647_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_647_inst_req_1;
      type_cast_647_inst_ack_1<= rack(0);
      type_cast_647_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_647_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call8_258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_648,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_355_index_1_rename
    process(R_indvar_354_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_354_resized;
      ov(13 downto 0) := iv;
      R_indvar_354_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_355_index_1_resize
    process(indvar_343) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_343;
      ov := iv(13 downto 0);
      R_indvar_354_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_355_root_address_inst
    process(array_obj_ref_355_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_355_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_355_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_492_addr_0
    process(ptr_deref_492_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_492_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_492_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_492_base_resize
    process(arrayidx_357) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_357;
      ov := iv(13 downto 0);
      ptr_deref_492_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_492_gather_scatter
    process(add61_490) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add61_490;
      ov(63 downto 0) := iv;
      ptr_deref_492_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_492_root_address_inst
    process(ptr_deref_492_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_492_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_492_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_293_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp126_292;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_293_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_293_branch_req_0,
          ack0 => if_stmt_293_branch_ack_0,
          ack1 => if_stmt_293_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_506_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond8_505;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_506_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_506_branch_req_0,
          ack0 => if_stmt_506_branch_ack_0,
          ack1 => if_stmt_506_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_499_inst
    process(indvar_343) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_343, type_cast_498_wire_constant, tmp_var);
      indvarx_xnext_500 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_285_inst
    process(mul13_280) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul13_280, type_cast_284_wire_constant, tmp_var);
      shr125x_xmask_286 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_291_inst
    process(shr125x_xmask_286) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr125x_xmask_286, type_cast_290_wire_constant, tmp_var);
      cmp126_292 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_504_inst
    process(indvarx_xnext_500, umax7_340) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_500, umax7_340, tmp_var);
      exitcond8_505 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_326_inst
    process(tmp4_321) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_321, type_cast_325_wire_constant, tmp_var);
      tmp5_327 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_652_inst
    process(conv118_644, conv116_640) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv118_644, conv116_640, tmp_var);
      mul119_653 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_657_inst
    process(mul119_653, conv121_648) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul119_653, conv121_648, tmp_var);
      mul122_658 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_274_inst
    process(conv10_266, conv_262) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv10_266, conv_262, tmp_var);
      mul_275 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_279_inst
    process(mul_275, conv12_270) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_275, conv12_270, tmp_var);
      mul13_280 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_311_inst
    process(tmp_303, tmp1_307) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_303, tmp1_307, tmp_var);
      tmp2_312 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_320_inst
    process(tmp2_312, tmp3_316) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_312, tmp3_316, tmp_var);
      tmp4_321 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_381_inst
    process(shl_370, conv25_377) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_370, conv25_377, tmp_var);
      add_382 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_399_inst
    process(shl27_388, conv30_395) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_388, conv30_395, tmp_var);
      add31_400 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_417_inst
    process(shl33_406, conv36_413) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl33_406, conv36_413, tmp_var);
      add37_418 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_435_inst
    process(shl39_424, conv42_431) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl39_424, conv42_431, tmp_var);
      add43_436 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_453_inst
    process(shl45_442, conv48_449) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_442, conv48_449, tmp_var);
      add49_454 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_471_inst
    process(shl51_460, conv54_467) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl51_460, conv54_467, tmp_var);
      add55_472 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_489_inst
    process(shl57_478, conv60_485) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl57_478, conv60_485, tmp_var);
      add61_490 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_369_inst
    process(conv21_364) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv21_364, type_cast_368_wire_constant, tmp_var);
      shl_370 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_387_inst
    process(add_382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_382, type_cast_386_wire_constant, tmp_var);
      shl27_388 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_405_inst
    process(add31_400) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add31_400, type_cast_404_wire_constant, tmp_var);
      shl33_406 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_423_inst
    process(add37_418) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add37_418, type_cast_422_wire_constant, tmp_var);
      shl39_424 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_441_inst
    process(add43_436) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add43_436, type_cast_440_wire_constant, tmp_var);
      shl45_442 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_459_inst
    process(add49_454) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add49_454, type_cast_458_wire_constant, tmp_var);
      shl51_460 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_477_inst
    process(add55_472) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add55_472, type_cast_476_wire_constant, tmp_var);
      shl57_478 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_631_inst
    process(conv110_627, conv67_523) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv110_627, conv67_523, tmp_var);
      sub_632 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_332_inst
    process(tmp5_327) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp5_327, type_cast_331_wire_constant, tmp_var);
      tmp6_333 <= tmp_var; --
    end process;
    -- shared split operator group (27) : array_obj_ref_355_index_offset 
    ApIntAdd_group_27: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_354_scaled;
      array_obj_ref_355_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_355_index_offset_req_0;
      array_obj_ref_355_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_355_index_offset_req_1;
      array_obj_ref_355_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_27_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_27_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- unary operator type_cast_521_inst
    process(call66_517) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call66_517, tmp_var);
      type_cast_521_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_625_inst
    process(call109_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call109_622, tmp_var);
      type_cast_625_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_492_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_492_store_0_req_0;
      ptr_deref_492_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_492_store_0_req_1;
      ptr_deref_492_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_492_word_address_0;
      data_in <= ptr_deref_492_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_complete_609_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_complete_609_inst_req_0;
      RPIPE_Block0_complete_609_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_complete_609_inst_req_1;
      RPIPE_Block0_complete_609_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call97_610 <= data_out(7 downto 0);
      Block0_complete_read_0_gI: SplitGuardInterface generic map(name => "Block0_complete_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_complete_read_0: InputPortRevised -- 
        generic map ( name => "Block0_complete_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_complete_pipe_read_req(0),
          oack => Block0_complete_pipe_read_ack(0),
          odata => Block0_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_complete_612_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_complete_612_inst_req_0;
      RPIPE_Block1_complete_612_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_complete_612_inst_req_1;
      RPIPE_Block1_complete_612_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call100_613 <= data_out(7 downto 0);
      Block1_complete_read_1_gI: SplitGuardInterface generic map(name => "Block1_complete_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_complete_read_1: InputPortRevised -- 
        generic map ( name => "Block1_complete_read_1", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_complete_pipe_read_req(0),
          oack => Block1_complete_pipe_read_ack(0),
          odata => Block1_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_complete_615_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_complete_615_inst_req_0;
      RPIPE_Block2_complete_615_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_complete_615_inst_req_1;
      RPIPE_Block2_complete_615_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call103_616 <= data_out(7 downto 0);
      Block2_complete_read_2_gI: SplitGuardInterface generic map(name => "Block2_complete_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_complete_read_2: InputPortRevised -- 
        generic map ( name => "Block2_complete_read_2", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_complete_pipe_read_req(0),
          oack => Block2_complete_pipe_read_ack(0),
          odata => Block2_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_complete_618_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_complete_618_inst_req_0;
      RPIPE_Block3_complete_618_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_complete_618_inst_req_1;
      RPIPE_Block3_complete_618_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call106_619 <= data_out(7 downto 0);
      Block3_complete_read_3_gI: SplitGuardInterface generic map(name => "Block3_complete_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_complete_read_3: InputPortRevised -- 
        generic map ( name => "Block3_complete_read_3", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_complete_pipe_read_req(0),
          oack => Block3_complete_pipe_read_ack(0),
          odata => Block3_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_zeropad_input_pipe_233_inst RPIPE_zeropad_input_pipe_236_inst RPIPE_zeropad_input_pipe_239_inst RPIPE_zeropad_input_pipe_242_inst RPIPE_zeropad_input_pipe_245_inst RPIPE_zeropad_input_pipe_248_inst RPIPE_zeropad_input_pipe_251_inst RPIPE_zeropad_input_pipe_254_inst RPIPE_zeropad_input_pipe_257_inst RPIPE_zeropad_input_pipe_359_inst RPIPE_zeropad_input_pipe_372_inst RPIPE_zeropad_input_pipe_390_inst RPIPE_zeropad_input_pipe_408_inst RPIPE_zeropad_input_pipe_426_inst RPIPE_zeropad_input_pipe_444_inst RPIPE_zeropad_input_pipe_462_inst RPIPE_zeropad_input_pipe_480_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(135 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 16 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 16 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 16 downto 0);
      signal guard_vector : std_logic_vector( 16 downto 0);
      constant outBUFs : IntegerArray(16 downto 0) := (16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(16 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false);
      constant guardBuffering: IntegerArray(16 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2);
      -- 
    begin -- 
      reqL_unguarded(16) <= RPIPE_zeropad_input_pipe_233_inst_req_0;
      reqL_unguarded(15) <= RPIPE_zeropad_input_pipe_236_inst_req_0;
      reqL_unguarded(14) <= RPIPE_zeropad_input_pipe_239_inst_req_0;
      reqL_unguarded(13) <= RPIPE_zeropad_input_pipe_242_inst_req_0;
      reqL_unguarded(12) <= RPIPE_zeropad_input_pipe_245_inst_req_0;
      reqL_unguarded(11) <= RPIPE_zeropad_input_pipe_248_inst_req_0;
      reqL_unguarded(10) <= RPIPE_zeropad_input_pipe_251_inst_req_0;
      reqL_unguarded(9) <= RPIPE_zeropad_input_pipe_254_inst_req_0;
      reqL_unguarded(8) <= RPIPE_zeropad_input_pipe_257_inst_req_0;
      reqL_unguarded(7) <= RPIPE_zeropad_input_pipe_359_inst_req_0;
      reqL_unguarded(6) <= RPIPE_zeropad_input_pipe_372_inst_req_0;
      reqL_unguarded(5) <= RPIPE_zeropad_input_pipe_390_inst_req_0;
      reqL_unguarded(4) <= RPIPE_zeropad_input_pipe_408_inst_req_0;
      reqL_unguarded(3) <= RPIPE_zeropad_input_pipe_426_inst_req_0;
      reqL_unguarded(2) <= RPIPE_zeropad_input_pipe_444_inst_req_0;
      reqL_unguarded(1) <= RPIPE_zeropad_input_pipe_462_inst_req_0;
      reqL_unguarded(0) <= RPIPE_zeropad_input_pipe_480_inst_req_0;
      RPIPE_zeropad_input_pipe_233_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_zeropad_input_pipe_236_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_zeropad_input_pipe_239_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_zeropad_input_pipe_242_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_zeropad_input_pipe_245_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_zeropad_input_pipe_248_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_zeropad_input_pipe_251_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_zeropad_input_pipe_254_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_zeropad_input_pipe_257_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_zeropad_input_pipe_359_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_zeropad_input_pipe_372_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_zeropad_input_pipe_390_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_zeropad_input_pipe_408_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_zeropad_input_pipe_426_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_zeropad_input_pipe_444_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_zeropad_input_pipe_462_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_zeropad_input_pipe_480_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(16) <= RPIPE_zeropad_input_pipe_233_inst_req_1;
      reqR_unguarded(15) <= RPIPE_zeropad_input_pipe_236_inst_req_1;
      reqR_unguarded(14) <= RPIPE_zeropad_input_pipe_239_inst_req_1;
      reqR_unguarded(13) <= RPIPE_zeropad_input_pipe_242_inst_req_1;
      reqR_unguarded(12) <= RPIPE_zeropad_input_pipe_245_inst_req_1;
      reqR_unguarded(11) <= RPIPE_zeropad_input_pipe_248_inst_req_1;
      reqR_unguarded(10) <= RPIPE_zeropad_input_pipe_251_inst_req_1;
      reqR_unguarded(9) <= RPIPE_zeropad_input_pipe_254_inst_req_1;
      reqR_unguarded(8) <= RPIPE_zeropad_input_pipe_257_inst_req_1;
      reqR_unguarded(7) <= RPIPE_zeropad_input_pipe_359_inst_req_1;
      reqR_unguarded(6) <= RPIPE_zeropad_input_pipe_372_inst_req_1;
      reqR_unguarded(5) <= RPIPE_zeropad_input_pipe_390_inst_req_1;
      reqR_unguarded(4) <= RPIPE_zeropad_input_pipe_408_inst_req_1;
      reqR_unguarded(3) <= RPIPE_zeropad_input_pipe_426_inst_req_1;
      reqR_unguarded(2) <= RPIPE_zeropad_input_pipe_444_inst_req_1;
      reqR_unguarded(1) <= RPIPE_zeropad_input_pipe_462_inst_req_1;
      reqR_unguarded(0) <= RPIPE_zeropad_input_pipe_480_inst_req_1;
      RPIPE_zeropad_input_pipe_233_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_zeropad_input_pipe_236_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_zeropad_input_pipe_239_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_zeropad_input_pipe_242_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_zeropad_input_pipe_245_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_zeropad_input_pipe_248_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_zeropad_input_pipe_251_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_zeropad_input_pipe_254_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_zeropad_input_pipe_257_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_zeropad_input_pipe_359_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_zeropad_input_pipe_372_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_zeropad_input_pipe_390_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_zeropad_input_pipe_408_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_zeropad_input_pipe_426_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_zeropad_input_pipe_444_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_zeropad_input_pipe_462_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_zeropad_input_pipe_480_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      call_234 <= data_out(135 downto 128);
      call1_237 <= data_out(127 downto 120);
      call2_240 <= data_out(119 downto 112);
      call3_243 <= data_out(111 downto 104);
      call4_246 <= data_out(103 downto 96);
      call5_249 <= data_out(95 downto 88);
      call6_252 <= data_out(87 downto 80);
      call7_255 <= data_out(79 downto 72);
      call8_258 <= data_out(71 downto 64);
      call20_360 <= data_out(63 downto 56);
      call23_373 <= data_out(55 downto 48);
      call28_391 <= data_out(47 downto 40);
      call34_409 <= data_out(39 downto 32);
      call40_427 <= data_out(31 downto 24);
      call46_445 <= data_out(23 downto 16);
      call52_463 <= data_out(15 downto 8);
      call58_481 <= data_out(7 downto 0);
      zeropad_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "zeropad_input_pipe_read_4_gI", nreqs => 17, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      zeropad_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "zeropad_input_pipe_read_4", data_width => 8,  num_reqs => 17,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => zeropad_input_pipe_pipe_read_req(0),
          oack => zeropad_input_pipe_pipe_read_ack(0),
          odata => zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_starting_524_inst WPIPE_Block0_starting_527_inst WPIPE_Block0_starting_530_inst WPIPE_Block0_starting_533_inst WPIPE_Block0_starting_536_inst WPIPE_Block0_starting_539_inst WPIPE_Block0_starting_542_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block0_starting_524_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_starting_527_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_starting_530_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_starting_533_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_starting_536_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_starting_539_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_starting_542_inst_req_0;
      WPIPE_Block0_starting_524_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_starting_527_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_starting_530_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_starting_533_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_starting_536_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_starting_539_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_starting_542_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block0_starting_524_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_starting_527_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_starting_530_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_starting_533_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_starting_536_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_starting_539_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_starting_542_inst_req_1;
      WPIPE_Block0_starting_524_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_starting_527_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_starting_530_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_starting_533_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_starting_536_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_starting_539_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_starting_542_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call2_240 & call3_243 & call4_246 & call6_252 & call7_255 & call8_258 & call5_249;
      Block0_starting_write_0_gI: SplitGuardInterface generic map(name => "Block0_starting_write_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_starting_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_starting_pipe_write_req(0),
          oack => Block0_starting_pipe_write_ack(0),
          odata => Block0_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_starting_545_inst WPIPE_Block1_starting_548_inst WPIPE_Block1_starting_551_inst WPIPE_Block1_starting_554_inst WPIPE_Block1_starting_557_inst WPIPE_Block1_starting_560_inst WPIPE_Block1_starting_563_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block1_starting_545_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_starting_548_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_starting_551_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_starting_554_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_starting_557_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_starting_560_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_starting_563_inst_req_0;
      WPIPE_Block1_starting_545_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_starting_548_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_starting_551_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_starting_554_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_starting_557_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_starting_560_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_starting_563_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block1_starting_545_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_starting_548_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_starting_551_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_starting_554_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_starting_557_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_starting_560_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_starting_563_inst_req_1;
      WPIPE_Block1_starting_545_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_starting_548_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_starting_551_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_starting_554_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_starting_557_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_starting_560_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_starting_563_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call2_240 & call3_243 & call4_246 & call6_252 & call7_255 & call8_258 & call5_249;
      Block1_starting_write_1_gI: SplitGuardInterface generic map(name => "Block1_starting_write_1_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_starting_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_starting_pipe_write_req(0),
          oack => Block1_starting_pipe_write_ack(0),
          odata => Block1_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_starting_566_inst WPIPE_Block2_starting_569_inst WPIPE_Block2_starting_572_inst WPIPE_Block2_starting_575_inst WPIPE_Block2_starting_578_inst WPIPE_Block2_starting_581_inst WPIPE_Block2_starting_584_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block2_starting_566_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_starting_569_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_starting_572_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_starting_575_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_starting_578_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_starting_581_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_starting_584_inst_req_0;
      WPIPE_Block2_starting_566_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_starting_569_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_starting_572_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_starting_575_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_starting_578_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_starting_581_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_starting_584_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block2_starting_566_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_starting_569_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_starting_572_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_starting_575_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_starting_578_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_starting_581_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_starting_584_inst_req_1;
      WPIPE_Block2_starting_566_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_starting_569_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_starting_572_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_starting_575_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_starting_578_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_starting_581_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_starting_584_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call2_240 & call3_243 & call4_246 & call6_252 & call7_255 & call8_258 & call5_249;
      Block2_starting_write_2_gI: SplitGuardInterface generic map(name => "Block2_starting_write_2_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_starting_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_starting_pipe_write_req(0),
          oack => Block2_starting_pipe_write_ack(0),
          odata => Block2_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_starting_587_inst WPIPE_Block3_starting_590_inst WPIPE_Block3_starting_593_inst WPIPE_Block3_starting_596_inst WPIPE_Block3_starting_599_inst WPIPE_Block3_starting_602_inst WPIPE_Block3_starting_605_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block3_starting_587_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_starting_590_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_starting_593_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_starting_596_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_starting_599_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_starting_602_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_starting_605_inst_req_0;
      WPIPE_Block3_starting_587_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_starting_590_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_starting_593_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_starting_596_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_starting_599_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_starting_602_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_starting_605_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block3_starting_587_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_starting_590_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_starting_593_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_starting_596_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_starting_599_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_starting_602_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_starting_605_inst_req_1;
      WPIPE_Block3_starting_587_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_starting_590_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_starting_593_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_starting_596_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_starting_599_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_starting_602_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_starting_605_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call2_240 & call3_243 & call4_246 & call6_252 & call7_255 & call8_258 & call5_249;
      Block3_starting_write_3_gI: SplitGuardInterface generic map(name => "Block3_starting_write_3_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_starting_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_starting_pipe_write_req(0),
          oack => Block3_starting_pipe_write_ack(0),
          odata => Block3_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_elapsed_time_pipe_633_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_633_inst_req_0;
      WPIPE_elapsed_time_pipe_633_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_633_inst_req_1;
      WPIPE_elapsed_time_pipe_633_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_632;
      elapsed_time_pipe_write_4_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_517_call call_stmt_622_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_517_call_req_0;
      reqL_unguarded(0) <= call_stmt_622_call_req_0;
      call_stmt_517_call_ack_0 <= ackL_unguarded(1);
      call_stmt_622_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_517_call_req_1;
      reqR_unguarded(0) <= call_stmt_622_call_req_1;
      call_stmt_517_call_ack_1 <= ackR_unguarded(1);
      call_stmt_622_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call66_517 <= data_out(127 downto 64);
      call109_622 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_660_call 
    sendOutput_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_660_call_req_0;
      call_stmt_660_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_660_call_req_1;
      call_stmt_660_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul122_658;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          dataR => sendOutput_call_data(31 downto 0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_A is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block0_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block0_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_A;
architecture zeropad3D_A_arch of zeropad3D_A is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_A_CP_1955_start: Boolean;
  signal zeropad3D_A_CP_1955_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1127_inst_ack_1 : boolean;
  signal type_cast_1110_inst_req_0 : boolean;
  signal ptr_deref_1030_load_0_req_0 : boolean;
  signal array_obj_ref_1050_index_offset_req_1 : boolean;
  signal type_cast_1044_inst_ack_0 : boolean;
  signal type_cast_1044_inst_ack_1 : boolean;
  signal ptr_deref_1030_load_0_req_1 : boolean;
  signal addr_of_1051_final_reg_req_0 : boolean;
  signal type_cast_1110_inst_req_1 : boolean;
  signal addr_of_1051_final_reg_ack_0 : boolean;
  signal ptr_deref_1054_store_0_req_0 : boolean;
  signal if_stmt_1134_branch_ack_0 : boolean;
  signal if_stmt_1077_branch_ack_0 : boolean;
  signal type_cast_1062_inst_req_1 : boolean;
  signal type_cast_1127_inst_req_1 : boolean;
  signal addr_of_1051_final_reg_ack_1 : boolean;
  signal if_stmt_1077_branch_req_0 : boolean;
  signal ptr_deref_1030_load_0_ack_1 : boolean;
  signal ptr_deref_1030_load_0_ack_0 : boolean;
  signal type_cast_1127_inst_req_0 : boolean;
  signal ptr_deref_1054_store_0_ack_0 : boolean;
  signal type_cast_1110_inst_ack_0 : boolean;
  signal type_cast_1044_inst_req_1 : boolean;
  signal if_stmt_1077_branch_ack_1 : boolean;
  signal addr_of_1051_final_reg_req_1 : boolean;
  signal WPIPE_Block0_complete_1164_inst_req_0 : boolean;
  signal array_obj_ref_1050_index_offset_req_0 : boolean;
  signal phi_stmt_797_req_1 : boolean;
  signal array_obj_ref_1050_index_offset_ack_1 : boolean;
  signal type_cast_801_inst_req_0 : boolean;
  signal type_cast_1127_inst_ack_0 : boolean;
  signal array_obj_ref_1050_index_offset_ack_0 : boolean;
  signal type_cast_1110_inst_ack_1 : boolean;
  signal if_stmt_1134_branch_req_0 : boolean;
  signal type_cast_801_inst_ack_0 : boolean;
  signal type_cast_1062_inst_ack_1 : boolean;
  signal WPIPE_Block0_complete_1164_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_668_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_671_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_674_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_674_inst_req_0 : boolean;
  signal ptr_deref_1054_store_0_ack_1 : boolean;
  signal RPIPE_Block0_starting_668_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_671_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_674_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_668_inst_req_0 : boolean;
  signal type_cast_1044_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_668_inst_ack_0 : boolean;
  signal type_cast_1062_inst_req_0 : boolean;
  signal type_cast_1062_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_671_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_671_inst_ack_1 : boolean;
  signal phi_stmt_812_req_0 : boolean;
  signal WPIPE_Block0_complete_1164_inst_req_1 : boolean;
  signal type_cast_1101_inst_req_0 : boolean;
  signal type_cast_1101_inst_ack_0 : boolean;
  signal WPIPE_Block0_complete_1164_inst_ack_1 : boolean;
  signal type_cast_1101_inst_req_1 : boolean;
  signal phi_stmt_805_req_0 : boolean;
  signal type_cast_1101_inst_ack_1 : boolean;
  signal ptr_deref_1054_store_0_req_1 : boolean;
  signal if_stmt_1134_branch_ack_1 : boolean;
  signal RPIPE_Block0_starting_674_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_677_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_677_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_677_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_677_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_680_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_680_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_680_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_680_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_683_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_683_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_683_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_683_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_686_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_686_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_686_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_686_inst_ack_1 : boolean;
  signal type_cast_691_inst_req_0 : boolean;
  signal type_cast_691_inst_ack_0 : boolean;
  signal type_cast_691_inst_req_1 : boolean;
  signal type_cast_691_inst_ack_1 : boolean;
  signal type_cast_695_inst_req_0 : boolean;
  signal type_cast_695_inst_ack_0 : boolean;
  signal type_cast_695_inst_req_1 : boolean;
  signal type_cast_695_inst_ack_1 : boolean;
  signal type_cast_699_inst_req_0 : boolean;
  signal type_cast_699_inst_ack_0 : boolean;
  signal type_cast_699_inst_req_1 : boolean;
  signal type_cast_699_inst_ack_1 : boolean;
  signal type_cast_703_inst_req_0 : boolean;
  signal type_cast_703_inst_ack_0 : boolean;
  signal type_cast_703_inst_req_1 : boolean;
  signal type_cast_703_inst_ack_1 : boolean;
  signal type_cast_712_inst_req_0 : boolean;
  signal type_cast_712_inst_ack_0 : boolean;
  signal type_cast_712_inst_req_1 : boolean;
  signal type_cast_712_inst_ack_1 : boolean;
  signal type_cast_716_inst_req_0 : boolean;
  signal type_cast_716_inst_ack_0 : boolean;
  signal type_cast_716_inst_req_1 : boolean;
  signal type_cast_716_inst_ack_1 : boolean;
  signal type_cast_752_inst_req_0 : boolean;
  signal type_cast_752_inst_ack_0 : boolean;
  signal type_cast_752_inst_req_1 : boolean;
  signal type_cast_752_inst_ack_1 : boolean;
  signal type_cast_823_inst_req_0 : boolean;
  signal type_cast_823_inst_ack_0 : boolean;
  signal type_cast_823_inst_req_1 : boolean;
  signal type_cast_823_inst_ack_1 : boolean;
  signal if_stmt_850_branch_req_0 : boolean;
  signal if_stmt_850_branch_ack_1 : boolean;
  signal if_stmt_850_branch_ack_0 : boolean;
  signal type_cast_860_inst_req_0 : boolean;
  signal type_cast_860_inst_ack_0 : boolean;
  signal type_cast_860_inst_req_1 : boolean;
  signal type_cast_860_inst_ack_1 : boolean;
  signal if_stmt_887_branch_req_0 : boolean;
  signal if_stmt_887_branch_ack_1 : boolean;
  signal if_stmt_887_branch_ack_0 : boolean;
  signal type_cast_897_inst_req_0 : boolean;
  signal type_cast_897_inst_ack_0 : boolean;
  signal type_cast_897_inst_req_1 : boolean;
  signal type_cast_897_inst_ack_1 : boolean;
  signal type_cast_902_inst_req_0 : boolean;
  signal type_cast_902_inst_ack_0 : boolean;
  signal type_cast_902_inst_req_1 : boolean;
  signal type_cast_902_inst_ack_1 : boolean;
  signal type_cast_936_inst_req_0 : boolean;
  signal type_cast_936_inst_ack_0 : boolean;
  signal type_cast_936_inst_req_1 : boolean;
  signal type_cast_936_inst_ack_1 : boolean;
  signal array_obj_ref_942_index_offset_req_0 : boolean;
  signal array_obj_ref_942_index_offset_ack_0 : boolean;
  signal array_obj_ref_942_index_offset_req_1 : boolean;
  signal array_obj_ref_942_index_offset_ack_1 : boolean;
  signal addr_of_943_final_reg_req_0 : boolean;
  signal addr_of_943_final_reg_ack_0 : boolean;
  signal addr_of_943_final_reg_req_1 : boolean;
  signal addr_of_943_final_reg_ack_1 : boolean;
  signal ptr_deref_946_store_0_req_0 : boolean;
  signal ptr_deref_946_store_0_ack_0 : boolean;
  signal ptr_deref_946_store_0_req_1 : boolean;
  signal ptr_deref_946_store_0_ack_1 : boolean;
  signal type_cast_955_inst_req_0 : boolean;
  signal type_cast_955_inst_ack_0 : boolean;
  signal type_cast_955_inst_req_1 : boolean;
  signal type_cast_955_inst_ack_1 : boolean;
  signal type_cast_1019_inst_req_0 : boolean;
  signal type_cast_1019_inst_ack_0 : boolean;
  signal type_cast_1019_inst_req_1 : boolean;
  signal type_cast_1019_inst_ack_1 : boolean;
  signal array_obj_ref_1025_index_offset_req_0 : boolean;
  signal array_obj_ref_1025_index_offset_ack_0 : boolean;
  signal array_obj_ref_1025_index_offset_req_1 : boolean;
  signal array_obj_ref_1025_index_offset_ack_1 : boolean;
  signal addr_of_1026_final_reg_req_0 : boolean;
  signal addr_of_1026_final_reg_ack_0 : boolean;
  signal addr_of_1026_final_reg_req_1 : boolean;
  signal addr_of_1026_final_reg_ack_1 : boolean;
  signal type_cast_801_inst_req_1 : boolean;
  signal type_cast_801_inst_ack_1 : boolean;
  signal phi_stmt_797_req_0 : boolean;
  signal type_cast_811_inst_req_0 : boolean;
  signal type_cast_811_inst_ack_0 : boolean;
  signal type_cast_811_inst_req_1 : boolean;
  signal type_cast_811_inst_ack_1 : boolean;
  signal phi_stmt_805_req_1 : boolean;
  signal type_cast_818_inst_req_0 : boolean;
  signal type_cast_818_inst_ack_0 : boolean;
  signal type_cast_818_inst_req_1 : boolean;
  signal type_cast_818_inst_ack_1 : boolean;
  signal phi_stmt_812_req_1 : boolean;
  signal phi_stmt_797_ack_0 : boolean;
  signal phi_stmt_805_ack_0 : boolean;
  signal phi_stmt_812_ack_0 : boolean;
  signal phi_stmt_1141_req_1 : boolean;
  signal type_cast_1153_inst_req_0 : boolean;
  signal type_cast_1153_inst_ack_0 : boolean;
  signal type_cast_1153_inst_req_1 : boolean;
  signal type_cast_1153_inst_ack_1 : boolean;
  signal phi_stmt_1148_req_1 : boolean;
  signal type_cast_1159_inst_req_0 : boolean;
  signal type_cast_1159_inst_ack_0 : boolean;
  signal type_cast_1159_inst_req_1 : boolean;
  signal type_cast_1159_inst_ack_1 : boolean;
  signal phi_stmt_1154_req_1 : boolean;
  signal type_cast_1144_inst_req_0 : boolean;
  signal type_cast_1144_inst_ack_0 : boolean;
  signal type_cast_1144_inst_req_1 : boolean;
  signal type_cast_1144_inst_ack_1 : boolean;
  signal phi_stmt_1141_req_0 : boolean;
  signal type_cast_1151_inst_req_0 : boolean;
  signal type_cast_1151_inst_ack_0 : boolean;
  signal type_cast_1151_inst_req_1 : boolean;
  signal type_cast_1151_inst_ack_1 : boolean;
  signal phi_stmt_1148_req_0 : boolean;
  signal type_cast_1157_inst_req_0 : boolean;
  signal type_cast_1157_inst_ack_0 : boolean;
  signal type_cast_1157_inst_req_1 : boolean;
  signal type_cast_1157_inst_ack_1 : boolean;
  signal phi_stmt_1154_req_0 : boolean;
  signal phi_stmt_1141_ack_0 : boolean;
  signal phi_stmt_1148_ack_0 : boolean;
  signal phi_stmt_1154_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_A_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_A_CP_1955_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_A_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_A_CP_1955_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_A_CP_1955_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_A_CP_1955_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_A_CP_1955: Block -- control-path 
    signal zeropad3D_A_CP_1955_elements: BooleanArray(130 downto 0);
    -- 
  begin -- 
    zeropad3D_A_CP_1955_elements(0) <= zeropad3D_A_CP_1955_start;
    zeropad3D_A_CP_1955_symbol <= zeropad3D_A_CP_1955_elements(86);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/$entry
      -- CP-element group 0: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687__entry__
      -- CP-element group 0: 	 branch_block_stmt_666/branch_block_stmt_666__entry__
      -- CP-element group 0: 	 branch_block_stmt_666/$entry
      -- CP-element group 0: 	 $entry
      -- 
    rr_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(0), ack => RPIPE_Block0_starting_668_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	130 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	94 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	97 
    -- CP-element group 1: 	98 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_666/merge_stmt_1140__exit__
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/SplitProtocol/Update/cr
      -- 
    rr_2828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(1), ack => type_cast_801_inst_req_0); -- 
    cr_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(1), ack => type_cast_801_inst_req_1); -- 
    rr_2851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(1), ack => type_cast_811_inst_req_0); -- 
    cr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(1), ack => type_cast_811_inst_req_1); -- 
    rr_2874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(1), ack => type_cast_818_inst_req_0); -- 
    cr_2879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(1), ack => type_cast_818_inst_req_1); -- 
    zeropad3D_A_CP_1955_elements(1) <= zeropad3D_A_CP_1955_elements(130);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_update_start_
      -- CP-element group 2: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_Sample/$exit
      -- 
    ra_2022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_668_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(2)); -- 
    cr_2026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(2), ack => RPIPE_Block0_starting_668_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_668_update_completed_
      -- 
    ca_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_668_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(3)); -- 
    rr_2035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(3), ack => RPIPE_Block0_starting_671_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_update_start_
      -- CP-element group 4: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_Update/$entry
      -- 
    ra_2036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_671_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(4)); -- 
    cr_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(4), ack => RPIPE_Block0_starting_671_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_671_Update/$exit
      -- 
    ca_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_671_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(5)); -- 
    rr_2049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(5), ack => RPIPE_Block0_starting_674_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_update_start_
      -- CP-element group 6: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_sample_completed_
      -- 
    ra_2050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_674_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(6)); -- 
    cr_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(6), ack => RPIPE_Block0_starting_674_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_674_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_Sample/rr
      -- 
    ca_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_674_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(7)); -- 
    rr_2063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(7), ack => RPIPE_Block0_starting_677_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_update_start_
      -- CP-element group 8: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_Update/cr
      -- 
    ra_2064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_677_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(8)); -- 
    cr_2068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(8), ack => RPIPE_Block0_starting_677_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_677_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_Sample/rr
      -- 
    ca_2069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_677_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(9)); -- 
    rr_2077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(9), ack => RPIPE_Block0_starting_680_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_update_start_
      -- CP-element group 10: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_Update/cr
      -- 
    ra_2078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_680_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(10)); -- 
    cr_2082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(10), ack => RPIPE_Block0_starting_680_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_680_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_Sample/rr
      -- 
    ca_2083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_680_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(11)); -- 
    rr_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(11), ack => RPIPE_Block0_starting_683_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_update_start_
      -- CP-element group 12: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_Update/cr
      -- 
    ra_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_683_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(12)); -- 
    cr_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(12), ack => RPIPE_Block0_starting_683_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_683_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_Sample/rr
      -- 
    ca_2097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_683_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(13)); -- 
    rr_2105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(13), ack => RPIPE_Block0_starting_686_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_update_start_
      -- CP-element group 14: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_Update/cr
      -- 
    ra_2106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_686_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(14)); -- 
    cr_2110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(14), ack => RPIPE_Block0_starting_686_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15:  members (49) 
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/$exit
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794__entry__
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687__exit__
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_669_to_assign_stmt_687/RPIPE_Block0_starting_686_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_update_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_update_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_update_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_update_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_update_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_update_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_update_start_
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_Update/cr
      -- 
    ca_2111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_686_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(15)); -- 
    rr_2122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_691_inst_req_0); -- 
    cr_2127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_691_inst_req_1); -- 
    rr_2136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_695_inst_req_0); -- 
    cr_2141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_695_inst_req_1); -- 
    rr_2150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_699_inst_req_0); -- 
    cr_2155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_699_inst_req_1); -- 
    rr_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_703_inst_req_0); -- 
    cr_2169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_703_inst_req_1); -- 
    rr_2178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_712_inst_req_0); -- 
    cr_2183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_712_inst_req_1); -- 
    rr_2192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_716_inst_req_0); -- 
    cr_2197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_716_inst_req_1); -- 
    rr_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_752_inst_req_0); -- 
    cr_2211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(15), ack => type_cast_752_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_Sample/ra
      -- 
    ra_2123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_691_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	30 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_691_Update/ca
      -- 
    ca_2128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_691_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_Sample/ra
      -- 
    ra_2137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_695_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	30 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_695_Update/ca
      -- 
    ca_2142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_695_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_Sample/ra
      -- 
    ra_2151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	30 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_699_Update/ca
      -- 
    ca_2156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_Sample/ra
      -- 
    ra_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_703_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	30 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_703_Update/ca
      -- 
    ca_2170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_703_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_Sample/ra
      -- 
    ra_2179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_712_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	30 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_712_Update/ca
      -- 
    ca_2184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_712_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_Sample/ra
      -- 
    ra_2193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_716_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_716_Update/ca
      -- 
    ca_2198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_716_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_Sample/ra
      -- 
    ra_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_752_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/type_cast_752_Update/ca
      -- 
    ca_2212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_752_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  place  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: 	19 
    -- CP-element group 30: 	21 
    -- CP-element group 30: 	23 
    -- CP-element group 30: 	25 
    -- CP-element group 30: 	27 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	87 
    -- CP-element group 30: 	88 
    -- CP-element group 30: 	89 
    -- CP-element group 30:  members (10) 
      -- CP-element group 30: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_805/$entry
      -- CP-element group 30: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_797/$entry
      -- CP-element group 30: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/$entry
      -- CP-element group 30: 	 branch_block_stmt_666/entry_whilex_xbody
      -- CP-element group 30: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794__exit__
      -- CP-element group 30: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/$entry
      -- CP-element group 30: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/$entry
      -- CP-element group 30: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 30: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_812/$entry
      -- CP-element group 30: 	 branch_block_stmt_666/assign_stmt_692_to_assign_stmt_794/$exit
      -- 
    zeropad3D_A_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(17) & zeropad3D_A_CP_1955_elements(19) & zeropad3D_A_CP_1955_elements(21) & zeropad3D_A_CP_1955_elements(23) & zeropad3D_A_CP_1955_elements(25) & zeropad3D_A_CP_1955_elements(27) & zeropad3D_A_CP_1955_elements(29);
      gj_zeropad3D_A_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	105 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_Sample/ra
      -- 
    ra_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_823_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(31)); -- 
    -- CP-element group 32:  branch  transition  place  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	105 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (13) 
      -- CP-element group 32: 	 branch_block_stmt_666/if_stmt_850__entry__
      -- CP-element group 32: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849__exit__
      -- CP-element group 32: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/$exit
      -- CP-element group 32: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_666/if_stmt_850_dead_link/$entry
      -- CP-element group 32: 	 branch_block_stmt_666/if_stmt_850_eval_test/$entry
      -- CP-element group 32: 	 branch_block_stmt_666/if_stmt_850_eval_test/$exit
      -- CP-element group 32: 	 branch_block_stmt_666/if_stmt_850_eval_test/branch_req
      -- CP-element group 32: 	 branch_block_stmt_666/R_orx_xcond_851_place
      -- CP-element group 32: 	 branch_block_stmt_666/if_stmt_850_if_link/$entry
      -- CP-element group 32: 	 branch_block_stmt_666/if_stmt_850_else_link/$entry
      -- 
    ca_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_823_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(32)); -- 
    branch_req_2237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(32), ack => if_stmt_850_branch_req_0); -- 
    -- CP-element group 33:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (18) 
      -- CP-element group 33: 	 branch_block_stmt_666/merge_stmt_856_PhiReqMerge
      -- CP-element group 33: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886__entry__
      -- CP-element group 33: 	 branch_block_stmt_666/merge_stmt_856__exit__
      -- CP-element group 33: 	 branch_block_stmt_666/if_stmt_850_if_link/$exit
      -- CP-element group 33: 	 branch_block_stmt_666/if_stmt_850_if_link/if_choice_transition
      -- CP-element group 33: 	 branch_block_stmt_666/whilex_xbody_lorx_xlhsx_xfalse54
      -- CP-element group 33: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/$entry
      -- CP-element group 33: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_update_start_
      -- CP-element group 33: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_666/whilex_xbody_lorx_xlhsx_xfalse54_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_666/whilex_xbody_lorx_xlhsx_xfalse54_PhiReq/$exit
      -- CP-element group 33: 	 branch_block_stmt_666/merge_stmt_856_PhiAck/$entry
      -- CP-element group 33: 	 branch_block_stmt_666/merge_stmt_856_PhiAck/$exit
      -- CP-element group 33: 	 branch_block_stmt_666/merge_stmt_856_PhiAck/dummy
      -- 
    if_choice_transition_2242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_850_branch_ack_1, ack => zeropad3D_A_CP_1955_elements(33)); -- 
    rr_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(33), ack => type_cast_860_inst_req_0); -- 
    cr_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(33), ack => type_cast_860_inst_req_1); -- 
    -- CP-element group 34:  transition  place  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	106 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_666/if_stmt_850_else_link/$exit
      -- CP-element group 34: 	 branch_block_stmt_666/if_stmt_850_else_link/else_choice_transition
      -- CP-element group 34: 	 branch_block_stmt_666/whilex_xbody_ifx_xthen
      -- CP-element group 34: 	 branch_block_stmt_666/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_666/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_850_branch_ack_0, ack => zeropad3D_A_CP_1955_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_Sample/ra
      -- 
    ra_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_860_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(35)); -- 
    -- CP-element group 36:  branch  transition  place  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (13) 
      -- CP-element group 36: 	 branch_block_stmt_666/if_stmt_887__entry__
      -- CP-element group 36: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886__exit__
      -- CP-element group 36: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/$exit
      -- CP-element group 36: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_666/assign_stmt_861_to_assign_stmt_886/type_cast_860_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_666/if_stmt_887_dead_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_666/if_stmt_887_eval_test/$entry
      -- CP-element group 36: 	 branch_block_stmt_666/if_stmt_887_eval_test/$exit
      -- CP-element group 36: 	 branch_block_stmt_666/if_stmt_887_eval_test/branch_req
      -- CP-element group 36: 	 branch_block_stmt_666/R_orx_xcond186_888_place
      -- CP-element group 36: 	 branch_block_stmt_666/if_stmt_887_if_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_666/if_stmt_887_else_link/$entry
      -- 
    ca_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_860_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(36)); -- 
    branch_req_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(36), ack => if_stmt_887_branch_req_0); -- 
    -- CP-element group 37:  fork  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	60 
    -- CP-element group 37: 	58 
    -- CP-element group 37: 	56 
    -- CP-element group 37: 	53 
    -- CP-element group 37: 	54 
    -- CP-element group 37: 	62 
    -- CP-element group 37: 	64 
    -- CP-element group 37: 	66 
    -- CP-element group 37: 	68 
    -- CP-element group 37: 	71 
    -- CP-element group 37:  members (46) 
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_final_index_sum_regn_Update/req
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/word_access_complete/word_0/cr
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Update/word_access_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_final_index_sum_regn_update_start
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_complete/req
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_update_start_
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/word_access_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_final_index_sum_regn_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/merge_stmt_951_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_update_start_
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056__entry__
      -- CP-element group 37: 	 branch_block_stmt_666/merge_stmt_951__exit__
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Update/word_access_complete/word_0/cr
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_update_start_
      -- CP-element group 37: 	 branch_block_stmt_666/if_stmt_887_if_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_666/if_stmt_887_if_link/if_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_666/lorx_xlhsx_xfalse54_ifx_xelse
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_update_start_
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_update_start_
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_update_start_
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_final_index_sum_regn_update_start
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_final_index_sum_regn_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_final_index_sum_regn_Update/req
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_complete/req
      -- CP-element group 37: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_update_start_
      -- CP-element group 37: 	 branch_block_stmt_666/lorx_xlhsx_xfalse54_ifx_xelse_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/lorx_xlhsx_xfalse54_ifx_xelse_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_666/merge_stmt_951_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_666/merge_stmt_951_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_666/merge_stmt_951_PhiAck/dummy
      -- 
    if_choice_transition_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_887_branch_ack_1, ack => zeropad3D_A_CP_1955_elements(37)); -- 
    req_2596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(37), ack => array_obj_ref_1050_index_offset_req_1); -- 
    cr_2546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(37), ack => ptr_deref_1030_load_0_req_1); -- 
    cr_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(37), ack => type_cast_1044_inst_req_1); -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(37), ack => addr_of_1051_final_reg_req_1); -- 
    cr_2661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(37), ack => ptr_deref_1054_store_0_req_1); -- 
    rr_2436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(37), ack => type_cast_955_inst_req_0); -- 
    cr_2441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(37), ack => type_cast_955_inst_req_1); -- 
    cr_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(37), ack => type_cast_1019_inst_req_1); -- 
    req_2486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(37), ack => array_obj_ref_1025_index_offset_req_1); -- 
    req_2501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(37), ack => addr_of_1026_final_reg_req_1); -- 
    -- CP-element group 38:  transition  place  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	106 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_666/if_stmt_887_else_link/$exit
      -- CP-element group 38: 	 branch_block_stmt_666/if_stmt_887_else_link/else_choice_transition
      -- CP-element group 38: 	 branch_block_stmt_666/lorx_xlhsx_xfalse54_ifx_xthen
      -- CP-element group 38: 	 branch_block_stmt_666/lorx_xlhsx_xfalse54_ifx_xthen_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_666/lorx_xlhsx_xfalse54_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_2282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_887_branch_ack_0, ack => zeropad3D_A_CP_1955_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	106 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_Sample/ra
      -- 
    ra_2296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_897_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	106 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_Update/ca
      -- 
    ca_2301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_897_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	106 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_Sample/ra
      -- 
    ra_2310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_902_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	106 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_Update/ca
      -- 
    ca_2315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_902_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_Sample/rr
      -- 
    rr_2323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(43), ack => type_cast_936_inst_req_0); -- 
    zeropad3D_A_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(40) & zeropad3D_A_CP_1955_elements(42);
      gj_zeropad3D_A_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_Sample/ra
      -- 
    ra_2324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_936_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	106 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_final_index_sum_regn_Sample/req
      -- 
    ca_2329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_936_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(45)); -- 
    req_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(45), ack => array_obj_ref_942_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	52 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_final_index_sum_regn_Sample/ack
      -- 
    ack_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_942_index_offset_ack_0, ack => zeropad3D_A_CP_1955_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	106 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_request/req
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_942_index_offset_ack_1, ack => zeropad3D_A_CP_1955_elements(47)); -- 
    req_2369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(47), ack => addr_of_943_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_request/ack
      -- 
    ack_2370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_943_final_reg_ack_0, ack => zeropad3D_A_CP_1955_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	106 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (28) 
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_word_addrgen/root_register_ack
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/ptr_deref_946_Split/$entry
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/ptr_deref_946_Split/$exit
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/ptr_deref_946_Split/split_req
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/ptr_deref_946_Split/split_ack
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/word_access_start/$entry
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/word_access_start/word_0/$entry
      -- CP-element group 49: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/word_access_start/word_0/rr
      -- 
    ack_2375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_943_final_reg_ack_1, ack => zeropad3D_A_CP_1955_elements(49)); -- 
    rr_2413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(49), ack => ptr_deref_946_store_0_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/word_access_start/$exit
      -- CP-element group 50: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Sample/word_access_start/word_0/ra
      -- 
    ra_2414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_946_store_0_ack_0, ack => zeropad3D_A_CP_1955_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	106 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Update/word_access_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Update/word_access_complete/word_0/ca
      -- 
    ca_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_946_store_0_ack_1, ack => zeropad3D_A_CP_1955_elements(51)); -- 
    -- CP-element group 52:  join  transition  place  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	46 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	107 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_666/ifx_xthen_ifx_xend
      -- CP-element group 52: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949__exit__
      -- CP-element group 52: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/$exit
      -- CP-element group 52: 	 branch_block_stmt_666/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_666/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(46) & zeropad3D_A_CP_1955_elements(51);
      gj_zeropad3D_A_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	37 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_Sample/ra
      -- 
    ra_2437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_955_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(53)); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	37 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	63 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_955_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_Sample/rr
      -- 
    ca_2442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_955_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(54)); -- 
    rr_2450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(54), ack => type_cast_1019_inst_req_0); -- 
    rr_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(54), ack => type_cast_1044_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_Sample/ra
      -- 
    ra_2451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1019_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	37 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (16) 
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1019_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_final_index_sum_regn_Sample/req
      -- 
    ca_2456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1019_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(56)); -- 
    req_2481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(56), ack => array_obj_ref_1025_index_offset_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	72 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_final_index_sum_regn_Sample/ack
      -- 
    ack_2482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1025_index_offset_ack_0, ack => zeropad3D_A_CP_1955_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	37 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1025_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_request/req
      -- 
    ack_2487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1025_index_offset_ack_1, ack => zeropad3D_A_CP_1955_elements(58)); -- 
    req_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(58), ack => addr_of_1026_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_request/ack
      -- 
    ack_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1026_final_reg_ack_0, ack => zeropad3D_A_CP_1955_elements(59)); -- 
    -- CP-element group 60:  join  fork  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	37 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (24) 
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Sample/word_access_start/word_0/rr
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_word_addrgen/root_register_ack
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Sample/word_access_start/$entry
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Sample/word_access_start/word_0/$entry
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1026_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_base_plus_offset/$entry
      -- 
    ack_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1026_final_reg_ack_1, ack => zeropad3D_A_CP_1955_elements(60)); -- 
    rr_2535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(60), ack => ptr_deref_1030_load_0_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Sample/word_access_start/$exit
      -- CP-element group 61: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Sample/word_access_start/word_0/ra
      -- CP-element group 61: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Sample/word_access_start/word_0/$exit
      -- CP-element group 61: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_sample_completed_
      -- 
    ra_2536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_load_0_ack_0, ack => zeropad3D_A_CP_1955_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	37 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	69 
    -- CP-element group 62:  members (9) 
      -- CP-element group 62: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/word_access_complete/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/word_access_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/word_access_complete/word_0/ca
      -- CP-element group 62: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/ptr_deref_1030_Merge/$exit
      -- CP-element group 62: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/ptr_deref_1030_Merge/$entry
      -- CP-element group 62: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/ptr_deref_1030_Merge/merge_req
      -- CP-element group 62: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_Update/ptr_deref_1030_Merge/merge_ack
      -- CP-element group 62: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1030_update_completed_
      -- 
    ca_2547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_load_0_ack_1, ack => zeropad3D_A_CP_1955_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	54 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_sample_completed_
      -- 
    ra_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1044_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	37 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (16) 
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_final_index_sum_regn_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_scale_1/scale_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_final_index_sum_regn_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_scale_1/$exit
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_scale_1/scale_rename_req
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_computed_1
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_resize_1/$entry
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_resize_1/$exit
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_resize_1/index_resize_ack
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_resize_1/index_resize_req
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_scale_1/$entry
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_resized_1
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_index_scaled_1
      -- CP-element group 64: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/type_cast_1044_update_completed_
      -- 
    ca_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1044_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(64)); -- 
    req_2591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(64), ack => array_obj_ref_1050_index_offset_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	72 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_final_index_sum_regn_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_final_index_sum_regn_sample_complete
      -- CP-element group 65: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_final_index_sum_regn_Sample/ack
      -- 
    ack_2592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1050_index_offset_ack_0, ack => zeropad3D_A_CP_1955_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	37 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (11) 
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_base_plus_offset/sum_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_root_address_calculated
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_request/req
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_request/$entry
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_base_plus_offset/sum_rename_req
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_base_plus_offset/$exit
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_base_plus_offset/$entry
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_final_index_sum_regn_Update/ack
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_final_index_sum_regn_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/array_obj_ref_1050_offset_calculated
      -- 
    ack_2597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1050_index_offset_ack_1, ack => zeropad3D_A_CP_1955_elements(66)); -- 
    req_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(66), ack => addr_of_1051_final_reg_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_request/$exit
      -- CP-element group 67: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_request/ack
      -- CP-element group 67: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_sample_completed_
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1051_final_reg_ack_0, ack => zeropad3D_A_CP_1955_elements(67)); -- 
    -- CP-element group 68:  fork  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	37 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (19) 
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_complete/$exit
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/addr_of_1051_complete/ack
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_base_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_word_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_base_addr_resize/$exit
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_base_address_resized
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_base_addr_resize/$entry
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_base_addr_resize/base_resize_req
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_base_addr_resize/base_resize_ack
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_word_addrgen/$entry
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_word_addrgen/$exit
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_word_addrgen/root_register_req
      -- CP-element group 68: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_word_addrgen/root_register_ack
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1051_final_reg_ack_1, ack => zeropad3D_A_CP_1955_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	62 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (9) 
      -- CP-element group 69: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/word_access_start/word_0/rr
      -- CP-element group 69: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/word_access_start/word_0/$entry
      -- CP-element group 69: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/ptr_deref_1054_Split/$entry
      -- CP-element group 69: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/ptr_deref_1054_Split/$exit
      -- CP-element group 69: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/word_access_start/$entry
      -- CP-element group 69: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/ptr_deref_1054_Split/split_req
      -- CP-element group 69: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/ptr_deref_1054_Split/split_ack
      -- CP-element group 69: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/$entry
      -- 
    rr_2650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(69), ack => ptr_deref_1054_store_0_req_0); -- 
    zeropad3D_A_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(62) & zeropad3D_A_CP_1955_elements(68);
      gj_zeropad3D_A_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/word_access_start/word_0/$exit
      -- CP-element group 70: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/word_access_start/word_0/ra
      -- CP-element group 70: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/word_access_start/$exit
      -- CP-element group 70: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Sample/$exit
      -- 
    ra_2651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1054_store_0_ack_0, ack => zeropad3D_A_CP_1955_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	37 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Update/word_access_complete/$exit
      -- CP-element group 71: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Update/word_access_complete/word_0/ca
      -- CP-element group 71: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_Update/word_access_complete/word_0/$exit
      -- CP-element group 71: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/ptr_deref_1054_update_completed_
      -- 
    ca_2662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1054_store_0_ack_1, ack => zeropad3D_A_CP_1955_elements(71)); -- 
    -- CP-element group 72:  join  transition  place  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	57 
    -- CP-element group 72: 	65 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	107 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_666/ifx_xelse_ifx_xend
      -- CP-element group 72: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056__exit__
      -- CP-element group 72: 	 branch_block_stmt_666/assign_stmt_956_to_assign_stmt_1056/$exit
      -- CP-element group 72: 	 branch_block_stmt_666/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_666/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(57) & zeropad3D_A_CP_1955_elements(65) & zeropad3D_A_CP_1955_elements(71);
      gj_zeropad3D_A_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	107 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_Sample/ra
      -- 
    ra_2674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1062_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	107 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_666/if_stmt_1077_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_666/if_stmt_1077_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_666/if_stmt_1077_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_666/if_stmt_1077_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_666/if_stmt_1077_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/$exit
      -- CP-element group 74: 	 branch_block_stmt_666/if_stmt_1077__entry__
      -- CP-element group 74: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076__exit__
      -- CP-element group 74: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_666/R_cmp139_1078_place
      -- CP-element group 74: 	 branch_block_stmt_666/if_stmt_1077_else_link/$entry
      -- 
    ca_2679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1062_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(74)); -- 
    branch_req_2687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(74), ack => if_stmt_1077_branch_req_0); -- 
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	116 
    -- CP-element group 75: 	117 
    -- CP-element group 75: 	119 
    -- CP-element group 75: 	120 
    -- CP-element group 75: 	122 
    -- CP-element group 75: 	123 
    -- CP-element group 75:  members (40) 
      -- CP-element group 75: 	 branch_block_stmt_666/if_stmt_1077_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xend_ifx_xthen141
      -- CP-element group 75: 	 branch_block_stmt_666/if_stmt_1077_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180
      -- CP-element group 75: 	 branch_block_stmt_666/assign_stmt_1089__exit__
      -- CP-element group 75: 	 branch_block_stmt_666/assign_stmt_1089__entry__
      -- CP-element group 75: 	 branch_block_stmt_666/merge_stmt_1083__exit__
      -- CP-element group 75: 	 branch_block_stmt_666/merge_stmt_1083_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_666/assign_stmt_1089/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/assign_stmt_1089/$exit
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xend_ifx_xthen141_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xend_ifx_xthen141_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_666/merge_stmt_1083_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/merge_stmt_1083_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_666/merge_stmt_1083_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/SplitProtocol/Update/cr
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/SplitProtocol/Update/cr
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1077_branch_ack_1, ack => zeropad3D_A_CP_1955_elements(75)); -- 
    rr_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(75), ack => type_cast_1144_inst_req_0); -- 
    cr_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(75), ack => type_cast_1144_inst_req_1); -- 
    rr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(75), ack => type_cast_1151_inst_req_0); -- 
    cr_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(75), ack => type_cast_1151_inst_req_1); -- 
    rr_3080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(75), ack => type_cast_1157_inst_req_0); -- 
    cr_3085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(75), ack => type_cast_1157_inst_req_1); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76: 	80 
    -- CP-element group 76: 	82 
    -- CP-element group 76:  members (24) 
      -- CP-element group 76: 	 branch_block_stmt_666/if_stmt_1077_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/$entry
      -- CP-element group 76: 	 branch_block_stmt_666/if_stmt_1077_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_666/ifx_xend_ifx_xelse146
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_666/merge_stmt_1091_PhiReqMerge
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133__entry__
      -- CP-element group 76: 	 branch_block_stmt_666/merge_stmt_1091__exit__
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_update_start_
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_update_start_
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_update_start_
      -- CP-element group 76: 	 branch_block_stmt_666/ifx_xend_ifx_xelse146_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_666/ifx_xend_ifx_xelse146_PhiReq/$exit
      -- CP-element group 76: 	 branch_block_stmt_666/merge_stmt_1091_PhiAck/$entry
      -- CP-element group 76: 	 branch_block_stmt_666/merge_stmt_1091_PhiAck/$exit
      -- CP-element group 76: 	 branch_block_stmt_666/merge_stmt_1091_PhiAck/dummy
      -- 
    else_choice_transition_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1077_branch_ack_0, ack => zeropad3D_A_CP_1955_elements(76)); -- 
    cr_2731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(76), ack => type_cast_1110_inst_req_1); -- 
    cr_2745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(76), ack => type_cast_1127_inst_req_1); -- 
    rr_2712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(76), ack => type_cast_1101_inst_req_0); -- 
    cr_2717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(76), ack => type_cast_1101_inst_req_1); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_Sample/ra
      -- 
    ra_2713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1101_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1101_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_sample_start_
      -- 
    ca_2718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1101_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(78)); -- 
    rr_2726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(78), ack => type_cast_1110_inst_req_0); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_sample_completed_
      -- 
    ra_2727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	76 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1110_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_Sample/$entry
      -- 
    ca_2732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(80)); -- 
    rr_2740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(80), ack => type_cast_1127_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_Sample/$exit
      -- 
    ra_2741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1127_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(81)); -- 
    -- CP-element group 82:  branch  transition  place  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	76 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (13) 
      -- CP-element group 82: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_666/if_stmt_1134_dead_link/$entry
      -- CP-element group 82: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_666/R_cmp172_1135_place
      -- CP-element group 82: 	 branch_block_stmt_666/if_stmt_1134_eval_test/$entry
      -- CP-element group 82: 	 branch_block_stmt_666/if_stmt_1134_eval_test/$exit
      -- CP-element group 82: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/$exit
      -- CP-element group 82: 	 branch_block_stmt_666/if_stmt_1134_eval_test/branch_req
      -- CP-element group 82: 	 branch_block_stmt_666/if_stmt_1134_else_link/$entry
      -- CP-element group 82: 	 branch_block_stmt_666/if_stmt_1134__entry__
      -- CP-element group 82: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133__exit__
      -- CP-element group 82: 	 branch_block_stmt_666/if_stmt_1134_if_link/$entry
      -- CP-element group 82: 	 branch_block_stmt_666/assign_stmt_1097_to_assign_stmt_1133/type_cast_1127_update_completed_
      -- 
    ca_2746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1127_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(82)); -- 
    branch_req_2754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(82), ack => if_stmt_1134_branch_req_0); -- 
    -- CP-element group 83:  transition  place  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (15) 
      -- CP-element group 83: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_Sample/req
      -- CP-element group 83: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_666/assign_stmt_1167__entry__
      -- CP-element group 83: 	 branch_block_stmt_666/merge_stmt_1162__exit__
      -- CP-element group 83: 	 branch_block_stmt_666/assign_stmt_1167/$entry
      -- CP-element group 83: 	 branch_block_stmt_666/ifx_xelse146_whilex_xend
      -- CP-element group 83: 	 branch_block_stmt_666/if_stmt_1134_if_link/$exit
      -- CP-element group 83: 	 branch_block_stmt_666/if_stmt_1134_if_link/if_choice_transition
      -- CP-element group 83: 	 branch_block_stmt_666/ifx_xelse146_whilex_xend_PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_666/ifx_xelse146_whilex_xend_PhiReq/$exit
      -- CP-element group 83: 	 branch_block_stmt_666/merge_stmt_1162_PhiReqMerge
      -- CP-element group 83: 	 branch_block_stmt_666/merge_stmt_1162_PhiAck/$entry
      -- CP-element group 83: 	 branch_block_stmt_666/merge_stmt_1162_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_666/merge_stmt_1162_PhiAck/dummy
      -- 
    if_choice_transition_2759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1134_branch_ack_1, ack => zeropad3D_A_CP_1955_elements(83)); -- 
    req_2776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(83), ack => WPIPE_Block0_complete_1164_inst_req_0); -- 
    -- CP-element group 84:  fork  transition  place  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	108 
    -- CP-element group 84: 	109 
    -- CP-element group 84: 	110 
    -- CP-element group 84: 	112 
    -- CP-element group 84: 	113 
    -- CP-element group 84:  members (22) 
      -- CP-element group 84: 	 branch_block_stmt_666/if_stmt_1134_else_link/else_choice_transition
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180
      -- CP-element group 84: 	 branch_block_stmt_666/if_stmt_1134_else_link/$exit
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1141/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/SplitProtocol/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/SplitProtocol/Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/SplitProtocol/Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/SplitProtocol/Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/SplitProtocol/Update/cr
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/SplitProtocol/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/SplitProtocol/Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/SplitProtocol/Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/SplitProtocol/Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1134_branch_ack_0, ack => zeropad3D_A_CP_1955_elements(84)); -- 
    rr_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(84), ack => type_cast_1153_inst_req_0); -- 
    cr_2990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(84), ack => type_cast_1153_inst_req_1); -- 
    rr_3008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(84), ack => type_cast_1159_inst_req_0); -- 
    cr_3013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(84), ack => type_cast_1159_inst_req_1); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_update_start_
      -- CP-element group 85: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_Sample/ack
      -- CP-element group 85: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_Update/req
      -- 
    ack_2777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_complete_1164_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(85)); -- 
    req_2781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(85), ack => WPIPE_Block0_complete_1164_inst_req_1); -- 
    -- CP-element group 86:  transition  place  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (16) 
      -- CP-element group 86: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_666/assign_stmt_1167/$exit
      -- CP-element group 86: 	 branch_block_stmt_666/merge_stmt_1169__exit__
      -- CP-element group 86: 	 branch_block_stmt_666/return__
      -- CP-element group 86: 	 branch_block_stmt_666/assign_stmt_1167__exit__
      -- CP-element group 86: 	 branch_block_stmt_666/branch_block_stmt_666__exit__
      -- CP-element group 86: 	 branch_block_stmt_666/$exit
      -- CP-element group 86: 	 $exit
      -- CP-element group 86: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_666/assign_stmt_1167/WPIPE_Block0_complete_1164_Update/ack
      -- CP-element group 86: 	 branch_block_stmt_666/return___PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_666/return___PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_666/merge_stmt_1169_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_666/merge_stmt_1169_PhiAck/$entry
      -- CP-element group 86: 	 branch_block_stmt_666/merge_stmt_1169_PhiAck/$exit
      -- CP-element group 86: 	 branch_block_stmt_666/merge_stmt_1169_PhiAck/dummy
      -- 
    ack_2782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_complete_1164_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(86)); -- 
    -- CP-element group 87:  transition  output  delay-element  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	30 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_797/$exit
      -- CP-element group 87: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_req
      -- CP-element group 87: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_804_konst_delay_trans
      -- CP-element group 87: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/$exit
      -- 
    phi_stmt_797_req_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_797_req_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(87), ack => phi_stmt_797_req_1); -- 
    -- Element group zeropad3D_A_CP_1955_elements(87) is a control-delay.
    cp_element_87_delay: control_delay_element  generic map(name => " 87_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_1955_elements(30), ack => zeropad3D_A_CP_1955_elements(87), clk => clk, reset =>reset);
    -- CP-element group 88:  transition  output  delay-element  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	30 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_805/$exit
      -- CP-element group 88: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_809_konst_delay_trans
      -- CP-element group 88: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_req
      -- 
    phi_stmt_805_req_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_805_req_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(88), ack => phi_stmt_805_req_0); -- 
    -- Element group zeropad3D_A_CP_1955_elements(88) is a control-delay.
    cp_element_88_delay: control_delay_element  generic map(name => " 88_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_1955_elements(30), ack => zeropad3D_A_CP_1955_elements(88), clk => clk, reset =>reset);
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	30 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_816_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_req
      -- CP-element group 89: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/phi_stmt_812/$exit
      -- 
    phi_stmt_812_req_2809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_812_req_2809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(89), ack => phi_stmt_812_req_0); -- 
    -- Element group zeropad3D_A_CP_1955_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_1955_elements(30), ack => zeropad3D_A_CP_1955_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  join  transition  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	101 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_666/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(87) & zeropad3D_A_CP_1955_elements(88) & zeropad3D_A_CP_1955_elements(89);
      gj_zeropad3D_A_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/SplitProtocol/Sample/ra
      -- 
    ra_2829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_801_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/SplitProtocol/Update/ca
      -- 
    ca_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_801_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	100 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/$exit
      -- CP-element group 93: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/$exit
      -- CP-element group 93: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_sources/type_cast_801/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_797/phi_stmt_797_req
      -- 
    phi_stmt_797_req_2835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_797_req_2835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(93), ack => phi_stmt_797_req_0); -- 
    zeropad3D_A_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(91) & zeropad3D_A_CP_1955_elements(92);
      gj_zeropad3D_A_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/SplitProtocol/Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/SplitProtocol/Sample/ra
      -- 
    ra_2852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_811_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/SplitProtocol/Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/SplitProtocol/Update/ca
      -- 
    ca_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_811_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/$exit
      -- CP-element group 96: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/$exit
      -- CP-element group 96: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_sources/type_cast_811/SplitProtocol/$exit
      -- CP-element group 96: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_805/phi_stmt_805_req
      -- 
    phi_stmt_805_req_2858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_805_req_2858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(96), ack => phi_stmt_805_req_1); -- 
    zeropad3D_A_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(94) & zeropad3D_A_CP_1955_elements(95);
      gj_zeropad3D_A_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	1 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/SplitProtocol/Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/SplitProtocol/Sample/ra
      -- 
    ra_2875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_818_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	1 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/SplitProtocol/Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/SplitProtocol/Update/ca
      -- 
    ca_2880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_818_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/$exit
      -- CP-element group 99: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/$exit
      -- CP-element group 99: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/$exit
      -- CP-element group 99: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_sources/type_cast_818/SplitProtocol/$exit
      -- CP-element group 99: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/phi_stmt_812/phi_stmt_812_req
      -- 
    phi_stmt_812_req_2881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_812_req_2881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(99), ack => phi_stmt_812_req_1); -- 
    zeropad3D_A_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(97) & zeropad3D_A_CP_1955_elements(98);
      gj_zeropad3D_A_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	93 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_666/ifx_xend180_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(93) & zeropad3D_A_CP_1955_elements(96) & zeropad3D_A_CP_1955_elements(99);
      gj_zeropad3D_A_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  merge  fork  transition  place  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	90 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101: 	103 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_666/merge_stmt_796_PhiReqMerge
      -- CP-element group 101: 	 branch_block_stmt_666/merge_stmt_796_PhiAck/$entry
      -- 
    zeropad3D_A_CP_1955_elements(101) <= OrReduce(zeropad3D_A_CP_1955_elements(90) & zeropad3D_A_CP_1955_elements(100));
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	105 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_666/merge_stmt_796_PhiAck/phi_stmt_797_ack
      -- 
    phi_stmt_797_ack_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_797_ack_0, ack => zeropad3D_A_CP_1955_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_666/merge_stmt_796_PhiAck/phi_stmt_805_ack
      -- 
    phi_stmt_805_ack_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_805_ack_0, ack => zeropad3D_A_CP_1955_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	101 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_666/merge_stmt_796_PhiAck/phi_stmt_812_ack
      -- 
    phi_stmt_812_ack_2888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_812_ack_0, ack => zeropad3D_A_CP_1955_elements(104)); -- 
    -- CP-element group 105:  join  fork  transition  place  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	102 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	31 
    -- CP-element group 105: 	32 
    -- CP-element group 105:  members (10) 
      -- CP-element group 105: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849__entry__
      -- CP-element group 105: 	 branch_block_stmt_666/merge_stmt_796__exit__
      -- CP-element group 105: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/$entry
      -- CP-element group 105: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_update_start_
      -- CP-element group 105: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_666/assign_stmt_824_to_assign_stmt_849/type_cast_823_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_666/merge_stmt_796_PhiAck/$exit
      -- 
    rr_2223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(105), ack => type_cast_823_inst_req_0); -- 
    cr_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(105), ack => type_cast_823_inst_req_1); -- 
    zeropad3D_A_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(102) & zeropad3D_A_CP_1955_elements(103) & zeropad3D_A_CP_1955_elements(104);
      gj_zeropad3D_A_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  merge  fork  transition  place  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	34 
    -- CP-element group 106: 	38 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	47 
    -- CP-element group 106: 	49 
    -- CP-element group 106: 	51 
    -- CP-element group 106: 	39 
    -- CP-element group 106: 	40 
    -- CP-element group 106: 	41 
    -- CP-element group 106: 	42 
    -- CP-element group 106: 	45 
    -- CP-element group 106:  members (33) 
      -- CP-element group 106: 	 branch_block_stmt_666/merge_stmt_893_PhiReqMerge
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949__entry__
      -- CP-element group 106: 	 branch_block_stmt_666/merge_stmt_893__exit__
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_update_start_
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_Sample/rr
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_897_Update/cr
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_update_start_
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_Sample/rr
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_902_Update/cr
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_update_start_
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/type_cast_936_Update/cr
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_update_start_
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_final_index_sum_regn_update_start
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_final_index_sum_regn_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/array_obj_ref_942_final_index_sum_regn_Update/req
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_complete/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/addr_of_943_complete/req
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_update_start_
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Update/word_access_complete/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Update/word_access_complete/word_0/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/assign_stmt_898_to_assign_stmt_949/ptr_deref_946_Update/word_access_complete/word_0/cr
      -- CP-element group 106: 	 branch_block_stmt_666/merge_stmt_893_PhiAck/$entry
      -- CP-element group 106: 	 branch_block_stmt_666/merge_stmt_893_PhiAck/$exit
      -- CP-element group 106: 	 branch_block_stmt_666/merge_stmt_893_PhiAck/dummy
      -- 
    rr_2295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(106), ack => type_cast_897_inst_req_0); -- 
    cr_2300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(106), ack => type_cast_897_inst_req_1); -- 
    rr_2309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(106), ack => type_cast_902_inst_req_0); -- 
    cr_2314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(106), ack => type_cast_902_inst_req_1); -- 
    cr_2328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(106), ack => type_cast_936_inst_req_1); -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(106), ack => array_obj_ref_942_index_offset_req_1); -- 
    req_2374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(106), ack => addr_of_943_final_reg_req_1); -- 
    cr_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(106), ack => ptr_deref_946_store_0_req_1); -- 
    zeropad3D_A_CP_1955_elements(106) <= OrReduce(zeropad3D_A_CP_1955_elements(34) & zeropad3D_A_CP_1955_elements(38));
    -- CP-element group 107:  merge  fork  transition  place  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	52 
    -- CP-element group 107: 	72 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	73 
    -- CP-element group 107: 	74 
    -- CP-element group 107:  members (13) 
      -- CP-element group 107: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_Update/cr
      -- CP-element group 107: 	 branch_block_stmt_666/merge_stmt_1058_PhiReqMerge
      -- CP-element group 107: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/$entry
      -- CP-element group 107: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076__entry__
      -- CP-element group 107: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_666/merge_stmt_1058__exit__
      -- CP-element group 107: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_update_start_
      -- CP-element group 107: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_666/assign_stmt_1063_to_assign_stmt_1076/type_cast_1062_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_666/merge_stmt_1058_PhiAck/$entry
      -- CP-element group 107: 	 branch_block_stmt_666/merge_stmt_1058_PhiAck/$exit
      -- CP-element group 107: 	 branch_block_stmt_666/merge_stmt_1058_PhiAck/dummy
      -- 
    cr_2678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(107), ack => type_cast_1062_inst_req_1); -- 
    rr_2673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(107), ack => type_cast_1062_inst_req_0); -- 
    zeropad3D_A_CP_1955_elements(107) <= OrReduce(zeropad3D_A_CP_1955_elements(52) & zeropad3D_A_CP_1955_elements(72));
    -- CP-element group 108:  transition  output  delay-element  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	84 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	115 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1141/$exit
      -- CP-element group 108: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1147_konst_delay_trans
      -- CP-element group 108: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_req
      -- 
    phi_stmt_1141_req_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1141_req_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(108), ack => phi_stmt_1141_req_1); -- 
    -- Element group zeropad3D_A_CP_1955_elements(108) is a control-delay.
    cp_element_108_delay: control_delay_element  generic map(name => " 108_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_1955_elements(84), ack => zeropad3D_A_CP_1955_elements(108), clk => clk, reset =>reset);
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	84 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/SplitProtocol/Sample/ra
      -- 
    ra_2986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1153_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	84 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/SplitProtocol/Update/ca
      -- 
    ca_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1153_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	115 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/$exit
      -- CP-element group 111: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/$exit
      -- CP-element group 111: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1153/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_req
      -- 
    phi_stmt_1148_req_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1148_req_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(111), ack => phi_stmt_1148_req_1); -- 
    zeropad3D_A_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(109) & zeropad3D_A_CP_1955_elements(110);
      gj_zeropad3D_A_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	84 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/SplitProtocol/Sample/ra
      -- 
    ra_3009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	84 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/SplitProtocol/Update/ca
      -- 
    ca_3014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/$exit
      -- CP-element group 114: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/$exit
      -- CP-element group 114: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1159/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_req
      -- 
    phi_stmt_1154_req_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1154_req_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(114), ack => phi_stmt_1154_req_1); -- 
    zeropad3D_A_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(112) & zeropad3D_A_CP_1955_elements(113);
      gj_zeropad3D_A_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	108 
    -- CP-element group 115: 	111 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	126 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_666/ifx_xelse146_ifx_xend180_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(108) & zeropad3D_A_CP_1955_elements(111) & zeropad3D_A_CP_1955_elements(114);
      gj_zeropad3D_A_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	75 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/SplitProtocol/Sample/ra
      -- 
    ra_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1144_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	75 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/SplitProtocol/Update/ca
      -- 
    ca_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1144_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	125 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/$exit
      -- CP-element group 118: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/$exit
      -- CP-element group 118: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_sources/type_cast_1144/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1141/phi_stmt_1141_req
      -- 
    phi_stmt_1141_req_3041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1141_req_3041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(118), ack => phi_stmt_1141_req_0); -- 
    zeropad3D_A_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(116) & zeropad3D_A_CP_1955_elements(117);
      gj_zeropad3D_A_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	75 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/SplitProtocol/Sample/ra
      -- 
    ra_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1151_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	75 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/SplitProtocol/Update/ca
      -- 
    ca_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1151_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	125 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/$exit
      -- CP-element group 121: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/$exit
      -- CP-element group 121: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_sources/type_cast_1151/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1148/phi_stmt_1148_req
      -- 
    phi_stmt_1148_req_3064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1148_req_3064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(121), ack => phi_stmt_1148_req_0); -- 
    zeropad3D_A_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(119) & zeropad3D_A_CP_1955_elements(120);
      gj_zeropad3D_A_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	75 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/SplitProtocol/Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/SplitProtocol/Sample/ra
      -- 
    ra_3081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1157_inst_ack_0, ack => zeropad3D_A_CP_1955_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	75 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/SplitProtocol/Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/SplitProtocol/Update/ca
      -- 
    ca_3086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1157_inst_ack_1, ack => zeropad3D_A_CP_1955_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/$exit
      -- CP-element group 124: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/$exit
      -- CP-element group 124: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/$exit
      -- CP-element group 124: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_sources/type_cast_1157/SplitProtocol/$exit
      -- CP-element group 124: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/phi_stmt_1154/phi_stmt_1154_req
      -- 
    phi_stmt_1154_req_3087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1154_req_3087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1955_elements(124), ack => phi_stmt_1154_req_0); -- 
    zeropad3D_A_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(122) & zeropad3D_A_CP_1955_elements(123);
      gj_zeropad3D_A_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	118 
    -- CP-element group 125: 	121 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_666/ifx_xthen141_ifx_xend180_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(118) & zeropad3D_A_CP_1955_elements(121) & zeropad3D_A_CP_1955_elements(124);
      gj_zeropad3D_A_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  merge  fork  transition  place  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	115 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126: 	129 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_666/merge_stmt_1140_PhiReqMerge
      -- CP-element group 126: 	 branch_block_stmt_666/merge_stmt_1140_PhiAck/$entry
      -- 
    zeropad3D_A_CP_1955_elements(126) <= OrReduce(zeropad3D_A_CP_1955_elements(115) & zeropad3D_A_CP_1955_elements(125));
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	130 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_666/merge_stmt_1140_PhiAck/phi_stmt_1141_ack
      -- 
    phi_stmt_1141_ack_3092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1141_ack_0, ack => zeropad3D_A_CP_1955_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_666/merge_stmt_1140_PhiAck/phi_stmt_1148_ack
      -- 
    phi_stmt_1148_ack_3093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1148_ack_0, ack => zeropad3D_A_CP_1955_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	126 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_666/merge_stmt_1140_PhiAck/phi_stmt_1154_ack
      -- 
    phi_stmt_1154_ack_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1154_ack_0, ack => zeropad3D_A_CP_1955_elements(129)); -- 
    -- CP-element group 130:  join  transition  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	127 
    -- CP-element group 130: 	128 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	1 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_666/merge_stmt_1140_PhiAck/$exit
      -- 
    zeropad3D_A_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1955_elements(127) & zeropad3D_A_CP_1955_elements(128) & zeropad3D_A_CP_1955_elements(129);
      gj_zeropad3D_A_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1955_elements(130), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1013_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1038_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_730_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_792_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_930_wire : std_logic_vector(31 downto 0);
    signal R_idxprom126_1024_resized : std_logic_vector(13 downto 0);
    signal R_idxprom126_1024_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom131_1049_resized : std_logic_vector(13 downto 0);
    signal R_idxprom131_1049_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_941_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_941_scaled : std_logic_vector(13 downto 0);
    signal add107_986 : std_logic_vector(31 downto 0);
    signal add117_1001 : std_logic_vector(31 downto 0);
    signal add123_1006 : std_logic_vector(31 downto 0);
    signal add136_1069 : std_logic_vector(31 downto 0);
    signal add144_1089 : std_logic_vector(15 downto 0);
    signal add155_749 : std_logic_vector(31 downto 0);
    signal add171_764 : std_logic_vector(31 downto 0);
    signal add69_774 : std_logic_vector(31 downto 0);
    signal add80_918 : std_logic_vector(31 downto 0);
    signal add86_923 : std_logic_vector(31 downto 0);
    signal add98_981 : std_logic_vector(31 downto 0);
    signal add_769 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1025_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1050_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1050_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1050_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1050_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1050_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1050_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_942_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_942_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_942_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_942_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_942_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_942_root_address : std_logic_vector(13 downto 0);
    signal arrayidx127_1027 : std_logic_vector(31 downto 0);
    signal arrayidx132_1052 : std_logic_vector(31 downto 0);
    signal arrayidx_944 : std_logic_vector(31 downto 0);
    signal call1_672 : std_logic_vector(7 downto 0);
    signal call2_675 : std_logic_vector(7 downto 0);
    signal call3_678 : std_logic_vector(7 downto 0);
    signal call4_681 : std_logic_vector(7 downto 0);
    signal call5_684 : std_logic_vector(7 downto 0);
    signal call6_687 : std_logic_vector(7 downto 0);
    signal call_669 : std_logic_vector(7 downto 0);
    signal cmp139_1076 : std_logic_vector(0 downto 0);
    signal cmp156_1107 : std_logic_vector(0 downto 0);
    signal cmp172_1133 : std_logic_vector(0 downto 0);
    signal cmp52_844 : std_logic_vector(0 downto 0);
    signal cmp59_868 : std_logic_vector(0 downto 0);
    signal cmp59x_xnot_874 : std_logic_vector(0 downto 0);
    signal cmp70_881 : std_logic_vector(0 downto 0);
    signal cmp_831 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_837 : std_logic_vector(0 downto 0);
    signal conv100_794 : std_logic_vector(31 downto 0);
    signal conv135_1063 : std_logic_vector(31 downto 0);
    signal conv149_1102 : std_logic_vector(31 downto 0);
    signal conv164_1128 : std_logic_vector(31 downto 0);
    signal conv166_753 : std_logic_vector(31 downto 0);
    signal conv27_692 : std_logic_vector(31 downto 0);
    signal conv29_696 : std_logic_vector(31 downto 0);
    signal conv33_700 : std_logic_vector(31 downto 0);
    signal conv35_704 : std_logic_vector(31 downto 0);
    signal conv42_824 : std_logic_vector(31 downto 0);
    signal conv44_713 : std_logic_vector(31 downto 0);
    signal conv56_861 : std_logic_vector(31 downto 0);
    signal conv74_898 : std_logic_vector(31 downto 0);
    signal conv76_717 : std_logic_vector(31 downto 0);
    signal conv78_903 : std_logic_vector(31 downto 0);
    signal conv82_732 : std_logic_vector(31 downto 0);
    signal conv90_956 : std_logic_vector(31 downto 0);
    signal div152_738 : std_logic_vector(31 downto 0);
    signal div167_759 : std_logic_vector(31 downto 0);
    signal idxprom126_1020 : std_logic_vector(63 downto 0);
    signal idxprom131_1045 : std_logic_vector(63 downto 0);
    signal idxprom_937 : std_logic_vector(63 downto 0);
    signal inc161_1111 : std_logic_vector(15 downto 0);
    signal inc161x_xix_x2_1116 : std_logic_vector(15 downto 0);
    signal inc_1097 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_1148 : std_logic_vector(15 downto 0);
    signal ix_x2_805 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_1154 : std_logic_vector(15 downto 0);
    signal jx_x1_812 : std_logic_vector(15 downto 0);
    signal jx_x2_1123 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_1141 : std_logic_vector(15 downto 0);
    signal kx_x1_797 : std_logic_vector(15 downto 0);
    signal mul106_976 : std_logic_vector(31 downto 0);
    signal mul116_991 : std_logic_vector(31 downto 0);
    signal mul122_996 : std_logic_vector(31 downto 0);
    signal mul36_709 : std_logic_vector(31 downto 0);
    signal mul79_908 : std_logic_vector(31 downto 0);
    signal mul85_913 : std_logic_vector(31 downto 0);
    signal mul97_966 : std_logic_vector(31 downto 0);
    signal mul_780 : std_logic_vector(31 downto 0);
    signal orx_xcond186_886 : std_logic_vector(0 downto 0);
    signal orx_xcond_849 : std_logic_vector(0 downto 0);
    signal ptr_deref_1030_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1030_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1030_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1030_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1030_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1054_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1054_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1054_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1054_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1054_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1054_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_946_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_946_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_946_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_946_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_946_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_946_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext185_723 : std_logic_vector(31 downto 0);
    signal sext_785 : std_logic_vector(31 downto 0);
    signal shl_744 : std_logic_vector(31 downto 0);
    signal shr125_1015 : std_logic_vector(31 downto 0);
    signal shr130_1040 : std_logic_vector(31 downto 0);
    signal shr_932 : std_logic_vector(31 downto 0);
    signal sub105_971 : std_logic_vector(31 downto 0);
    signal sub_961 : std_logic_vector(31 downto 0);
    signal tmp128_1031 : std_logic_vector(63 downto 0);
    signal type_cast_1009_wire : std_logic_vector(31 downto 0);
    signal type_cast_1012_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1018_wire : std_logic_vector(63 downto 0);
    signal type_cast_1034_wire : std_logic_vector(31 downto 0);
    signal type_cast_1037_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1043_wire : std_logic_vector(63 downto 0);
    signal type_cast_1061_wire : std_logic_vector(31 downto 0);
    signal type_cast_1067_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1072_wire : std_logic_vector(31 downto 0);
    signal type_cast_1074_wire : std_logic_vector(31 downto 0);
    signal type_cast_1087_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1095_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1100_wire : std_logic_vector(31 downto 0);
    signal type_cast_1120_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1126_wire : std_logic_vector(31 downto 0);
    signal type_cast_1144_wire : std_logic_vector(15 downto 0);
    signal type_cast_1147_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1151_wire : std_logic_vector(15 downto 0);
    signal type_cast_1153_wire : std_logic_vector(15 downto 0);
    signal type_cast_1157_wire : std_logic_vector(15 downto 0);
    signal type_cast_1159_wire : std_logic_vector(15 downto 0);
    signal type_cast_1166_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_721_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_726_wire : std_logic_vector(31 downto 0);
    signal type_cast_729_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_736_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_742_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_757_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_778_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_788_wire : std_logic_vector(31 downto 0);
    signal type_cast_791_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_801_wire : std_logic_vector(15 downto 0);
    signal type_cast_804_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_809_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_811_wire : std_logic_vector(15 downto 0);
    signal type_cast_816_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_818_wire : std_logic_vector(15 downto 0);
    signal type_cast_822_wire : std_logic_vector(31 downto 0);
    signal type_cast_827_wire : std_logic_vector(31 downto 0);
    signal type_cast_829_wire : std_logic_vector(31 downto 0);
    signal type_cast_835_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_840_wire : std_logic_vector(31 downto 0);
    signal type_cast_842_wire : std_logic_vector(31 downto 0);
    signal type_cast_859_wire : std_logic_vector(31 downto 0);
    signal type_cast_864_wire : std_logic_vector(31 downto 0);
    signal type_cast_866_wire : std_logic_vector(31 downto 0);
    signal type_cast_872_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_877_wire : std_logic_vector(31 downto 0);
    signal type_cast_879_wire : std_logic_vector(31 downto 0);
    signal type_cast_896_wire : std_logic_vector(31 downto 0);
    signal type_cast_901_wire : std_logic_vector(31 downto 0);
    signal type_cast_926_wire : std_logic_vector(31 downto 0);
    signal type_cast_929_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_935_wire : std_logic_vector(63 downto 0);
    signal type_cast_948_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_954_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1025_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1025_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1025_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1025_resized_base_address <= "00000000000000";
    array_obj_ref_1050_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1050_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1050_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1050_resized_base_address <= "00000000000000";
    array_obj_ref_942_constant_part_of_offset <= "00000000000000";
    array_obj_ref_942_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_942_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_942_resized_base_address <= "00000000000000";
    ptr_deref_1030_word_offset_0 <= "00000000000000";
    ptr_deref_1054_word_offset_0 <= "00000000000000";
    ptr_deref_946_word_offset_0 <= "00000000000000";
    type_cast_1012_wire_constant <= "00000000000000000000000000000010";
    type_cast_1037_wire_constant <= "00000000000000000000000000000010";
    type_cast_1067_wire_constant <= "00000000000000000000000000000100";
    type_cast_1087_wire_constant <= "0000000000000100";
    type_cast_1095_wire_constant <= "0000000000000001";
    type_cast_1120_wire_constant <= "0000000000000000";
    type_cast_1147_wire_constant <= "0000000000000000";
    type_cast_1166_wire_constant <= "00000001";
    type_cast_721_wire_constant <= "00000000000000000000000000010000";
    type_cast_729_wire_constant <= "00000000000000000000000000010000";
    type_cast_736_wire_constant <= "00000000000000000000000000000001";
    type_cast_742_wire_constant <= "00000000000000000000000000000001";
    type_cast_757_wire_constant <= "00000000000000000000000000000001";
    type_cast_778_wire_constant <= "00000000000000000000000000010000";
    type_cast_791_wire_constant <= "00000000000000000000000000010000";
    type_cast_804_wire_constant <= "0000000000000000";
    type_cast_809_wire_constant <= "0000000000000000";
    type_cast_816_wire_constant <= "0000000000000000";
    type_cast_835_wire_constant <= "1";
    type_cast_872_wire_constant <= "1";
    type_cast_929_wire_constant <= "00000000000000000000000000000010";
    type_cast_948_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1141: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1144_wire & type_cast_1147_wire_constant;
      req <= phi_stmt_1141_req_0 & phi_stmt_1141_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1141",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1141_ack_0,
          idata => idata,
          odata => kx_x0x_xph_1141,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1141
    phi_stmt_1148: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1151_wire & type_cast_1153_wire;
      req <= phi_stmt_1148_req_0 & phi_stmt_1148_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1148",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1148_ack_0,
          idata => idata,
          odata => ix_x1x_xph_1148,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1148
    phi_stmt_1154: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1157_wire & type_cast_1159_wire;
      req <= phi_stmt_1154_req_0 & phi_stmt_1154_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1154",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1154_ack_0,
          idata => idata,
          odata => jx_x0x_xph_1154,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1154
    phi_stmt_797: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_801_wire & type_cast_804_wire_constant;
      req <= phi_stmt_797_req_0 & phi_stmt_797_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_797",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_797_ack_0,
          idata => idata,
          odata => kx_x1_797,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_797
    phi_stmt_805: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_809_wire_constant & type_cast_811_wire;
      req <= phi_stmt_805_req_0 & phi_stmt_805_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_805",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_805_ack_0,
          idata => idata,
          odata => ix_x2_805,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_805
    phi_stmt_812: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_816_wire_constant & type_cast_818_wire;
      req <= phi_stmt_812_req_0 & phi_stmt_812_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_812",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_812_ack_0,
          idata => idata,
          odata => jx_x1_812,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_812
    -- flow-through select operator MUX_1122_inst
    jx_x2_1123 <= type_cast_1120_wire_constant when (cmp156_1107(0) /=  '0') else inc_1097;
    addr_of_1026_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1026_final_reg_req_0;
      addr_of_1026_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1026_final_reg_req_1;
      addr_of_1026_final_reg_ack_1<= rack(0);
      addr_of_1026_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1026_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1025_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx127_1027,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1051_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1051_final_reg_req_0;
      addr_of_1051_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1051_final_reg_req_1;
      addr_of_1051_final_reg_ack_1<= rack(0);
      addr_of_1051_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1051_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1050_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx132_1052,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_943_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_943_final_reg_req_0;
      addr_of_943_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_943_final_reg_req_1;
      addr_of_943_final_reg_ack_1<= rack(0);
      addr_of_943_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_943_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_942_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_944,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1009_inst
    process(add107_986) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add107_986(31 downto 0);
      type_cast_1009_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1014_inst
    process(ASHR_i32_i32_1013_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1013_wire(31 downto 0);
      shr125_1015 <= tmp_var; -- 
    end process;
    type_cast_1019_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1019_inst_req_0;
      type_cast_1019_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1019_inst_req_1;
      type_cast_1019_inst_ack_1<= rack(0);
      type_cast_1019_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1019_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1018_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom126_1020,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1034_inst
    process(add123_1006) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add123_1006(31 downto 0);
      type_cast_1034_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1039_inst
    process(ASHR_i32_i32_1038_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1038_wire(31 downto 0);
      shr130_1040 <= tmp_var; -- 
    end process;
    type_cast_1044_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1044_inst_req_0;
      type_cast_1044_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1044_inst_req_1;
      type_cast_1044_inst_ack_1<= rack(0);
      type_cast_1044_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1044_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1043_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom131_1045,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1062_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1062_inst_req_0;
      type_cast_1062_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1062_inst_req_1;
      type_cast_1062_inst_ack_1<= rack(0);
      type_cast_1062_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1062_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1061_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_1063,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1072_inst
    process(add136_1069) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add136_1069(31 downto 0);
      type_cast_1072_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1074_inst
    process(conv27_692) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv27_692(31 downto 0);
      type_cast_1074_wire <= tmp_var; -- 
    end process;
    type_cast_1101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1101_inst_req_0;
      type_cast_1101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1101_inst_req_1;
      type_cast_1101_inst_ack_1<= rack(0);
      type_cast_1101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1100_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_1102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1110_inst_req_0;
      type_cast_1110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1110_inst_req_1;
      type_cast_1110_inst_ack_1<= rack(0);
      type_cast_1110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp156_1107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc161_1111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1127_inst_req_0;
      type_cast_1127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1127_inst_req_1;
      type_cast_1127_inst_ack_1<= rack(0);
      type_cast_1127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1126_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv164_1128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1144_inst_req_0;
      type_cast_1144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1144_inst_req_1;
      type_cast_1144_inst_ack_1<= rack(0);
      type_cast_1144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add144_1089,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1144_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1151_inst_req_0;
      type_cast_1151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1151_inst_req_1;
      type_cast_1151_inst_ack_1<= rack(0);
      type_cast_1151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_805,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1151_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1153_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1153_inst_req_0;
      type_cast_1153_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1153_inst_req_1;
      type_cast_1153_inst_ack_1<= rack(0);
      type_cast_1153_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1153_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc161x_xix_x2_1116,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1153_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1157_inst_req_0;
      type_cast_1157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1157_inst_req_1;
      type_cast_1157_inst_ack_1<= rack(0);
      type_cast_1157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_812,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1157_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1159_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1159_inst_req_0;
      type_cast_1159_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1159_inst_req_1;
      type_cast_1159_inst_ack_1<= rack(0);
      type_cast_1159_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1159_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_1123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1159_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_691_inst_req_0;
      type_cast_691_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_691_inst_req_1;
      type_cast_691_inst_ack_1<= rack(0);
      type_cast_691_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_691_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_675,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_692,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_695_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_695_inst_req_0;
      type_cast_695_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_695_inst_req_1;
      type_cast_695_inst_ack_1<= rack(0);
      type_cast_695_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_695_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_672,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_696,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_699_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_699_inst_req_0;
      type_cast_699_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_699_inst_req_1;
      type_cast_699_inst_ack_1<= rack(0);
      type_cast_699_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_699_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_703_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_703_inst_req_0;
      type_cast_703_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_703_inst_req_1;
      type_cast_703_inst_ack_1<= rack(0);
      type_cast_703_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_703_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_681,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_704,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_712_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_712_inst_req_0;
      type_cast_712_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_712_inst_req_1;
      type_cast_712_inst_ack_1<= rack(0);
      type_cast_712_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_712_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_687,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_713,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_716_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_716_inst_req_0;
      type_cast_716_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_716_inst_req_1;
      type_cast_716_inst_ack_1<= rack(0);
      type_cast_716_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_716_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_717,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_726_inst
    process(sext185_723) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext185_723(31 downto 0);
      type_cast_726_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_731_inst
    process(ASHR_i32_i32_730_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_730_wire(31 downto 0);
      conv82_732 <= tmp_var; -- 
    end process;
    type_cast_752_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_752_inst_req_0;
      type_cast_752_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_752_inst_req_1;
      type_cast_752_inst_ack_1<= rack(0);
      type_cast_752_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_752_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_669,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv166_753,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_788_inst
    process(sext_785) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_785(31 downto 0);
      type_cast_788_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_793_inst
    process(ASHR_i32_i32_792_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_792_wire(31 downto 0);
      conv100_794 <= tmp_var; -- 
    end process;
    type_cast_801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_801_inst_req_0;
      type_cast_801_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_801_inst_req_1;
      type_cast_801_inst_ack_1<= rack(0);
      type_cast_801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_1141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_801_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_811_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_811_inst_req_0;
      type_cast_811_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_811_inst_req_1;
      type_cast_811_inst_ack_1<= rack(0);
      type_cast_811_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_811_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_1148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_811_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_818_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_818_inst_req_0;
      type_cast_818_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_818_inst_req_1;
      type_cast_818_inst_ack_1<= rack(0);
      type_cast_818_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_818_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_1154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_818_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_823_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_823_inst_req_0;
      type_cast_823_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_823_inst_req_1;
      type_cast_823_inst_ack_1<= rack(0);
      type_cast_823_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_823_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_822_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_824,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_827_inst
    process(conv42_824) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv42_824(31 downto 0);
      type_cast_827_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_829_inst
    process(conv44_713) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv44_713(31 downto 0);
      type_cast_829_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_840_inst
    process(conv42_824) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv42_824(31 downto 0);
      type_cast_840_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_842_inst
    process(add_769) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_769(31 downto 0);
      type_cast_842_wire <= tmp_var; -- 
    end process;
    type_cast_860_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_860_inst_req_0;
      type_cast_860_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_860_inst_req_1;
      type_cast_860_inst_ack_1<= rack(0);
      type_cast_860_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_860_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_859_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_861,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_864_inst
    process(conv56_861) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv56_861(31 downto 0);
      type_cast_864_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_866_inst
    process(conv44_713) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv44_713(31 downto 0);
      type_cast_866_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_877_inst
    process(conv56_861) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv56_861(31 downto 0);
      type_cast_877_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_879_inst
    process(add69_774) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add69_774(31 downto 0);
      type_cast_879_wire <= tmp_var; -- 
    end process;
    type_cast_897_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_897_inst_req_0;
      type_cast_897_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_897_inst_req_1;
      type_cast_897_inst_ack_1<= rack(0);
      type_cast_897_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_897_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_896_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_898,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_902_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_902_inst_req_0;
      type_cast_902_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_902_inst_req_1;
      type_cast_902_inst_ack_1<= rack(0);
      type_cast_902_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_902_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_901_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_903,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_926_inst
    process(add86_923) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add86_923(31 downto 0);
      type_cast_926_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_931_inst
    process(ASHR_i32_i32_930_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_930_wire(31 downto 0);
      shr_932 <= tmp_var; -- 
    end process;
    type_cast_936_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_936_inst_req_0;
      type_cast_936_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_936_inst_req_1;
      type_cast_936_inst_ack_1<= rack(0);
      type_cast_936_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_936_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_935_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_937,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_955_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_955_inst_req_0;
      type_cast_955_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_955_inst_req_1;
      type_cast_955_inst_ack_1<= rack(0);
      type_cast_955_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_955_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_954_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_956,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1025_index_1_rename
    process(R_idxprom126_1024_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom126_1024_resized;
      ov(13 downto 0) := iv;
      R_idxprom126_1024_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1025_index_1_resize
    process(idxprom126_1020) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom126_1020;
      ov := iv(13 downto 0);
      R_idxprom126_1024_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1025_root_address_inst
    process(array_obj_ref_1025_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1025_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1025_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1050_index_1_rename
    process(R_idxprom131_1049_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom131_1049_resized;
      ov(13 downto 0) := iv;
      R_idxprom131_1049_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1050_index_1_resize
    process(idxprom131_1045) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom131_1045;
      ov := iv(13 downto 0);
      R_idxprom131_1049_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1050_root_address_inst
    process(array_obj_ref_1050_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1050_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1050_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_942_index_1_rename
    process(R_idxprom_941_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_941_resized;
      ov(13 downto 0) := iv;
      R_idxprom_941_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_942_index_1_resize
    process(idxprom_937) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_937;
      ov := iv(13 downto 0);
      R_idxprom_941_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_942_root_address_inst
    process(array_obj_ref_942_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_942_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_942_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1030_addr_0
    process(ptr_deref_1030_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1030_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1030_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1030_base_resize
    process(arrayidx127_1027) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx127_1027;
      ov := iv(13 downto 0);
      ptr_deref_1030_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1030_gather_scatter
    process(ptr_deref_1030_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1030_data_0;
      ov(63 downto 0) := iv;
      tmp128_1031 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1030_root_address_inst
    process(ptr_deref_1030_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1030_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1030_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1054_addr_0
    process(ptr_deref_1054_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1054_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1054_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1054_base_resize
    process(arrayidx132_1052) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx132_1052;
      ov := iv(13 downto 0);
      ptr_deref_1054_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1054_gather_scatter
    process(tmp128_1031) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp128_1031;
      ov(63 downto 0) := iv;
      ptr_deref_1054_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1054_root_address_inst
    process(ptr_deref_1054_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1054_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1054_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_946_addr_0
    process(ptr_deref_946_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_946_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_946_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_946_base_resize
    process(arrayidx_944) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_944;
      ov := iv(13 downto 0);
      ptr_deref_946_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_946_gather_scatter
    process(type_cast_948_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_948_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_946_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_946_root_address_inst
    process(ptr_deref_946_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_946_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_946_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1077_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp139_1076;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1077_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1077_branch_req_0,
          ack0 => if_stmt_1077_branch_ack_0,
          ack1 => if_stmt_1077_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1134_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp172_1133;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1134_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1134_branch_req_0,
          ack0 => if_stmt_1134_branch_ack_0,
          ack1 => if_stmt_1134_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_850_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_849;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_850_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_850_branch_req_0,
          ack0 => if_stmt_850_branch_ack_0,
          ack1 => if_stmt_850_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_887_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond186_886;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_887_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_887_branch_req_0,
          ack0 => if_stmt_887_branch_ack_0,
          ack1 => if_stmt_887_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1088_inst
    process(kx_x1_797) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_797, type_cast_1087_wire_constant, tmp_var);
      add144_1089 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1096_inst
    process(jx_x1_812) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_812, type_cast_1095_wire_constant, tmp_var);
      inc_1097 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1115_inst
    process(inc161_1111, ix_x2_805) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc161_1111, ix_x2_805, tmp_var);
      inc161x_xix_x2_1116 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1000_inst
    process(mul122_996, conv90_956) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul122_996, conv90_956, tmp_var);
      add117_1001 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1005_inst
    process(add117_1001, mul116_991) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add117_1001, mul116_991, tmp_var);
      add123_1006 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1068_inst
    process(conv135_1063) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv135_1063, type_cast_1067_wire_constant, tmp_var);
      add136_1069 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_748_inst
    process(shl_744, div152_738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_744, div152_738, tmp_var);
      add155_749 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_763_inst
    process(shl_744, div167_759) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_744, div167_759, tmp_var);
      add171_764 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_768_inst
    process(conv44_713, div167_759) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv44_713, div167_759, tmp_var);
      add_769 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_773_inst
    process(conv44_713, div152_738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv44_713, div152_738, tmp_var);
      add69_774 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_917_inst
    process(mul85_913, conv74_898) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul85_913, conv74_898, tmp_var);
      add80_918 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_922_inst
    process(add80_918, mul79_908) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add80_918, mul79_908, tmp_var);
      add86_923 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_980_inst
    process(mul106_976, conv90_956) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul106_976, conv90_956, tmp_var);
      add98_981 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_985_inst
    process(add98_981, mul97_966) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add98_981, mul97_966, tmp_var);
      add107_986 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_848_inst
    process(cmpx_xnot_837, cmp52_844) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_837, cmp52_844, tmp_var);
      orx_xcond_849 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_885_inst
    process(cmp59x_xnot_874, cmp70_881) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp59x_xnot_874, cmp70_881, tmp_var);
      orx_xcond186_886 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1013_inst
    process(type_cast_1009_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1009_wire, type_cast_1012_wire_constant, tmp_var);
      ASHR_i32_i32_1013_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1038_inst
    process(type_cast_1034_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1034_wire, type_cast_1037_wire_constant, tmp_var);
      ASHR_i32_i32_1038_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_730_inst
    process(type_cast_726_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_726_wire, type_cast_729_wire_constant, tmp_var);
      ASHR_i32_i32_730_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_792_inst
    process(type_cast_788_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_788_wire, type_cast_791_wire_constant, tmp_var);
      ASHR_i32_i32_792_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_930_inst
    process(type_cast_926_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_926_wire, type_cast_929_wire_constant, tmp_var);
      ASHR_i32_i32_930_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1106_inst
    process(conv149_1102, add155_749) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv149_1102, add155_749, tmp_var);
      cmp156_1107 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1132_inst
    process(conv164_1128, add171_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv164_1128, add171_764, tmp_var);
      cmp172_1133 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_737_inst
    process(conv29_696) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv29_696, type_cast_736_wire_constant, tmp_var);
      div152_738 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_758_inst
    process(conv166_753) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv166_753, type_cast_757_wire_constant, tmp_var);
      div167_759 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_708_inst
    process(conv33_700, conv35_704) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv33_700, conv35_704, tmp_var);
      mul36_709 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_784_inst
    process(mul_780, conv27_692) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_780, conv27_692, tmp_var);
      sext_785 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_907_inst
    process(conv78_903, conv76_717) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv78_903, conv76_717, tmp_var);
      mul79_908 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_912_inst
    process(conv42_824, conv82_732) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv42_824, conv82_732, tmp_var);
      mul85_913 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_965_inst
    process(sub_961, conv27_692) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_961, conv27_692, tmp_var);
      mul97_966 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_975_inst
    process(sub105_971, conv100_794) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub105_971, conv100_794, tmp_var);
      mul106_976 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_990_inst
    process(conv56_861, conv76_717) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv56_861, conv76_717, tmp_var);
      mul116_991 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_995_inst
    process(conv42_824, conv82_732) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv42_824, conv82_732, tmp_var);
      mul122_996 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_722_inst
    process(mul36_709) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul36_709, type_cast_721_wire_constant, tmp_var);
      sext185_723 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_743_inst
    process(conv44_713) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_713, type_cast_742_wire_constant, tmp_var);
      shl_744 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_779_inst
    process(conv29_696) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_696, type_cast_778_wire_constant, tmp_var);
      mul_780 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1075_inst
    process(type_cast_1072_wire, type_cast_1074_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1072_wire, type_cast_1074_wire, tmp_var);
      cmp139_1076 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_830_inst
    process(type_cast_827_wire, type_cast_829_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_827_wire, type_cast_829_wire, tmp_var);
      cmp_831 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_843_inst
    process(type_cast_840_wire, type_cast_842_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_840_wire, type_cast_842_wire, tmp_var);
      cmp52_844 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_867_inst
    process(type_cast_864_wire, type_cast_866_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_864_wire, type_cast_866_wire, tmp_var);
      cmp59_868 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_880_inst
    process(type_cast_877_wire, type_cast_879_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_877_wire, type_cast_879_wire, tmp_var);
      cmp70_881 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_960_inst
    process(conv56_861, conv44_713) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv56_861, conv44_713, tmp_var);
      sub_961 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_970_inst
    process(conv42_824, conv44_713) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv42_824, conv44_713, tmp_var);
      sub105_971 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_836_inst
    process(cmp_831) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_831, type_cast_835_wire_constant, tmp_var);
      cmpx_xnot_837 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_873_inst
    process(cmp59_868) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp59_868, type_cast_872_wire_constant, tmp_var);
      cmp59x_xnot_874 <= tmp_var; --
    end process;
    -- shared split operator group (45) : array_obj_ref_1025_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom126_1024_scaled;
      array_obj_ref_1025_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1025_index_offset_req_0;
      array_obj_ref_1025_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1025_index_offset_req_1;
      array_obj_ref_1025_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : array_obj_ref_1050_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom131_1049_scaled;
      array_obj_ref_1050_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1050_index_offset_req_0;
      array_obj_ref_1050_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1050_index_offset_req_1;
      array_obj_ref_1050_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_942_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_941_scaled;
      array_obj_ref_942_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_942_index_offset_req_0;
      array_obj_ref_942_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_942_index_offset_req_1;
      array_obj_ref_942_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- unary operator type_cast_1018_inst
    process(shr125_1015) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr125_1015, tmp_var);
      type_cast_1018_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1043_inst
    process(shr130_1040) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr130_1040, tmp_var);
      type_cast_1043_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1061_inst
    process(kx_x1_797) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_797, tmp_var);
      type_cast_1061_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1100_inst
    process(inc_1097) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1097, tmp_var);
      type_cast_1100_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1126_inst
    process(inc161x_xix_x2_1116) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc161x_xix_x2_1116, tmp_var);
      type_cast_1126_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_822_inst
    process(ix_x2_805) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_805, tmp_var);
      type_cast_822_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_859_inst
    process(jx_x1_812) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_812, tmp_var);
      type_cast_859_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_896_inst
    process(kx_x1_797) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_797, tmp_var);
      type_cast_896_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_901_inst
    process(jx_x1_812) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_812, tmp_var);
      type_cast_901_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_935_inst
    process(shr_932) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_932, tmp_var);
      type_cast_935_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_954_inst
    process(kx_x1_797) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_797, tmp_var);
      type_cast_954_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1030_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1030_load_0_req_0;
      ptr_deref_1030_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1030_load_0_req_1;
      ptr_deref_1030_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1030_word_address_0;
      ptr_deref_1030_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_946_store_0 ptr_deref_1054_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_946_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1054_store_0_req_0;
      ptr_deref_946_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1054_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_946_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1054_store_0_req_1;
      ptr_deref_946_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1054_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_946_word_address_0 & ptr_deref_1054_word_address_0;
      data_in <= ptr_deref_946_data_0 & ptr_deref_1054_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_starting_674_inst RPIPE_Block0_starting_677_inst RPIPE_Block0_starting_680_inst RPIPE_Block0_starting_683_inst RPIPE_Block0_starting_686_inst RPIPE_Block0_starting_671_inst RPIPE_Block0_starting_668_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block0_starting_674_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_starting_677_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_starting_680_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_starting_683_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_starting_686_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_starting_671_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_starting_668_inst_req_0;
      RPIPE_Block0_starting_674_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_starting_677_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_starting_680_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_starting_683_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_starting_686_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_starting_671_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_starting_668_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block0_starting_674_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_starting_677_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_starting_680_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_starting_683_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_starting_686_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_starting_671_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_starting_668_inst_req_1;
      RPIPE_Block0_starting_674_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_starting_677_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_starting_680_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_starting_683_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_starting_686_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_starting_671_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_starting_668_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call2_675 <= data_out(55 downto 48);
      call3_678 <= data_out(47 downto 40);
      call4_681 <= data_out(39 downto 32);
      call5_684 <= data_out(31 downto 24);
      call6_687 <= data_out(23 downto 16);
      call1_672 <= data_out(15 downto 8);
      call_669 <= data_out(7 downto 0);
      Block0_starting_read_0_gI: SplitGuardInterface generic map(name => "Block0_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block0_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_starting_pipe_read_req(0),
          oack => Block0_starting_pipe_read_ack(0),
          odata => Block0_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_complete_1164_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_complete_1164_inst_req_0;
      WPIPE_Block0_complete_1164_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_complete_1164_inst_req_1;
      WPIPE_Block0_complete_1164_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1166_wire_constant;
      Block0_complete_write_0_gI: SplitGuardInterface generic map(name => "Block0_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_complete_pipe_write_req(0),
          oack => Block0_complete_pipe_write_ack(0),
          odata => Block0_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_A_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_B is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block1_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block1_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_B;
architecture zeropad3D_B_arch of zeropad3D_B is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_B_CP_3111_start: Boolean;
  signal zeropad3D_B_CP_3111_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1216_inst_ack_1 : boolean;
  signal type_cast_1369_inst_ack_0 : boolean;
  signal type_cast_1216_inst_req_1 : boolean;
  signal type_cast_1332_inst_ack_1 : boolean;
  signal if_stmt_1396_branch_ack_1 : boolean;
  signal type_cast_1216_inst_ack_0 : boolean;
  signal type_cast_1220_inst_ack_0 : boolean;
  signal type_cast_1332_inst_ack_0 : boolean;
  signal type_cast_1406_inst_ack_1 : boolean;
  signal type_cast_1332_inst_req_0 : boolean;
  signal type_cast_1406_inst_req_0 : boolean;
  signal type_cast_1369_inst_req_1 : boolean;
  signal if_stmt_1396_branch_ack_0 : boolean;
  signal type_cast_1233_inst_req_1 : boolean;
  signal type_cast_1369_inst_req_0 : boolean;
  signal type_cast_1233_inst_ack_1 : boolean;
  signal type_cast_1233_inst_ack_0 : boolean;
  signal if_stmt_1359_branch_ack_1 : boolean;
  signal type_cast_1445_inst_req_1 : boolean;
  signal type_cast_1445_inst_ack_0 : boolean;
  signal if_stmt_1359_branch_ack_0 : boolean;
  signal type_cast_1445_inst_ack_1 : boolean;
  signal type_cast_1229_inst_ack_0 : boolean;
  signal type_cast_1411_inst_req_0 : boolean;
  signal type_cast_1216_inst_req_0 : boolean;
  signal type_cast_1220_inst_req_0 : boolean;
  signal type_cast_1411_inst_ack_0 : boolean;
  signal type_cast_1263_inst_req_0 : boolean;
  signal type_cast_1229_inst_req_0 : boolean;
  signal type_cast_1332_inst_req_1 : boolean;
  signal type_cast_1411_inst_req_1 : boolean;
  signal type_cast_1369_inst_ack_1 : boolean;
  signal type_cast_1411_inst_ack_1 : boolean;
  signal type_cast_1263_inst_ack_0 : boolean;
  signal type_cast_1406_inst_ack_0 : boolean;
  signal type_cast_1233_inst_req_0 : boolean;
  signal type_cast_1229_inst_req_1 : boolean;
  signal type_cast_1263_inst_req_1 : boolean;
  signal type_cast_1406_inst_req_1 : boolean;
  signal type_cast_1445_inst_req_0 : boolean;
  signal if_stmt_1396_branch_req_0 : boolean;
  signal type_cast_1220_inst_req_1 : boolean;
  signal type_cast_1263_inst_ack_1 : boolean;
  signal type_cast_1220_inst_ack_1 : boolean;
  signal if_stmt_1359_branch_req_0 : boolean;
  signal array_obj_ref_1451_index_offset_req_1 : boolean;
  signal array_obj_ref_1451_index_offset_ack_1 : boolean;
  signal array_obj_ref_1451_index_offset_req_0 : boolean;
  signal array_obj_ref_1451_index_offset_ack_0 : boolean;
  signal type_cast_1229_inst_ack_1 : boolean;
  signal RPIPE_Block1_starting_1175_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1175_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1175_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1175_inst_ack_1 : boolean;
  signal RPIPE_Block1_starting_1178_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1178_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1178_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1178_inst_ack_1 : boolean;
  signal RPIPE_Block1_starting_1181_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1181_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1181_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1181_inst_ack_1 : boolean;
  signal RPIPE_Block1_starting_1184_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1184_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1184_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1184_inst_ack_1 : boolean;
  signal RPIPE_Block1_starting_1187_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1187_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1187_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1187_inst_ack_1 : boolean;
  signal RPIPE_Block1_starting_1190_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1190_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1190_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1190_inst_ack_1 : boolean;
  signal RPIPE_Block1_starting_1193_inst_req_0 : boolean;
  signal RPIPE_Block1_starting_1193_inst_ack_0 : boolean;
  signal RPIPE_Block1_starting_1193_inst_req_1 : boolean;
  signal RPIPE_Block1_starting_1193_inst_ack_1 : boolean;
  signal type_cast_1198_inst_req_0 : boolean;
  signal type_cast_1198_inst_ack_0 : boolean;
  signal type_cast_1198_inst_req_1 : boolean;
  signal type_cast_1198_inst_ack_1 : boolean;
  signal type_cast_1208_inst_req_0 : boolean;
  signal type_cast_1208_inst_ack_0 : boolean;
  signal type_cast_1208_inst_req_1 : boolean;
  signal type_cast_1208_inst_ack_1 : boolean;
  signal type_cast_1212_inst_req_0 : boolean;
  signal type_cast_1212_inst_ack_0 : boolean;
  signal type_cast_1212_inst_req_1 : boolean;
  signal type_cast_1212_inst_ack_1 : boolean;
  signal addr_of_1452_final_reg_req_0 : boolean;
  signal addr_of_1452_final_reg_ack_0 : boolean;
  signal addr_of_1452_final_reg_req_1 : boolean;
  signal addr_of_1452_final_reg_ack_1 : boolean;
  signal ptr_deref_1455_store_0_req_0 : boolean;
  signal ptr_deref_1455_store_0_ack_0 : boolean;
  signal ptr_deref_1455_store_0_req_1 : boolean;
  signal ptr_deref_1455_store_0_ack_1 : boolean;
  signal type_cast_1464_inst_req_0 : boolean;
  signal type_cast_1464_inst_ack_0 : boolean;
  signal type_cast_1464_inst_req_1 : boolean;
  signal type_cast_1464_inst_ack_1 : boolean;
  signal type_cast_1528_inst_req_0 : boolean;
  signal type_cast_1528_inst_ack_0 : boolean;
  signal type_cast_1528_inst_req_1 : boolean;
  signal type_cast_1528_inst_ack_1 : boolean;
  signal array_obj_ref_1534_index_offset_req_0 : boolean;
  signal array_obj_ref_1534_index_offset_ack_0 : boolean;
  signal array_obj_ref_1534_index_offset_req_1 : boolean;
  signal array_obj_ref_1534_index_offset_ack_1 : boolean;
  signal addr_of_1535_final_reg_req_0 : boolean;
  signal addr_of_1535_final_reg_ack_0 : boolean;
  signal addr_of_1535_final_reg_req_1 : boolean;
  signal addr_of_1535_final_reg_ack_1 : boolean;
  signal ptr_deref_1539_load_0_req_0 : boolean;
  signal ptr_deref_1539_load_0_ack_0 : boolean;
  signal ptr_deref_1539_load_0_req_1 : boolean;
  signal ptr_deref_1539_load_0_ack_1 : boolean;
  signal type_cast_1553_inst_req_0 : boolean;
  signal type_cast_1553_inst_ack_0 : boolean;
  signal type_cast_1553_inst_req_1 : boolean;
  signal type_cast_1553_inst_ack_1 : boolean;
  signal array_obj_ref_1559_index_offset_req_0 : boolean;
  signal array_obj_ref_1559_index_offset_ack_0 : boolean;
  signal array_obj_ref_1559_index_offset_req_1 : boolean;
  signal array_obj_ref_1559_index_offset_ack_1 : boolean;
  signal addr_of_1560_final_reg_req_0 : boolean;
  signal addr_of_1560_final_reg_ack_0 : boolean;
  signal addr_of_1560_final_reg_req_1 : boolean;
  signal addr_of_1560_final_reg_ack_1 : boolean;
  signal ptr_deref_1563_store_0_req_0 : boolean;
  signal ptr_deref_1563_store_0_ack_0 : boolean;
  signal ptr_deref_1563_store_0_req_1 : boolean;
  signal ptr_deref_1563_store_0_ack_1 : boolean;
  signal type_cast_1571_inst_req_0 : boolean;
  signal type_cast_1571_inst_ack_0 : boolean;
  signal type_cast_1571_inst_req_1 : boolean;
  signal type_cast_1571_inst_ack_1 : boolean;
  signal if_stmt_1586_branch_req_0 : boolean;
  signal if_stmt_1586_branch_ack_1 : boolean;
  signal if_stmt_1586_branch_ack_0 : boolean;
  signal type_cast_1610_inst_req_0 : boolean;
  signal type_cast_1610_inst_ack_0 : boolean;
  signal type_cast_1610_inst_req_1 : boolean;
  signal type_cast_1610_inst_ack_1 : boolean;
  signal type_cast_1619_inst_req_0 : boolean;
  signal type_cast_1619_inst_ack_0 : boolean;
  signal type_cast_1619_inst_req_1 : boolean;
  signal type_cast_1619_inst_ack_1 : boolean;
  signal type_cast_1635_inst_req_0 : boolean;
  signal type_cast_1635_inst_ack_0 : boolean;
  signal type_cast_1635_inst_req_1 : boolean;
  signal type_cast_1635_inst_ack_1 : boolean;
  signal if_stmt_1642_branch_req_0 : boolean;
  signal if_stmt_1642_branch_ack_1 : boolean;
  signal if_stmt_1642_branch_ack_0 : boolean;
  signal WPIPE_Block1_complete_1672_inst_req_0 : boolean;
  signal WPIPE_Block1_complete_1672_inst_ack_0 : boolean;
  signal WPIPE_Block1_complete_1672_inst_req_1 : boolean;
  signal WPIPE_Block1_complete_1672_inst_ack_1 : boolean;
  signal type_cast_1325_inst_req_0 : boolean;
  signal type_cast_1325_inst_ack_0 : boolean;
  signal type_cast_1325_inst_req_1 : boolean;
  signal type_cast_1325_inst_ack_1 : boolean;
  signal phi_stmt_1322_req_0 : boolean;
  signal phi_stmt_1308_req_0 : boolean;
  signal phi_stmt_1315_req_1 : boolean;
  signal type_cast_1327_inst_req_0 : boolean;
  signal type_cast_1327_inst_ack_0 : boolean;
  signal type_cast_1327_inst_req_1 : boolean;
  signal type_cast_1327_inst_ack_1 : boolean;
  signal phi_stmt_1322_req_1 : boolean;
  signal type_cast_1314_inst_req_0 : boolean;
  signal type_cast_1314_inst_ack_0 : boolean;
  signal type_cast_1314_inst_req_1 : boolean;
  signal type_cast_1314_inst_ack_1 : boolean;
  signal phi_stmt_1308_req_1 : boolean;
  signal type_cast_1318_inst_req_0 : boolean;
  signal type_cast_1318_inst_ack_0 : boolean;
  signal type_cast_1318_inst_req_1 : boolean;
  signal type_cast_1318_inst_ack_1 : boolean;
  signal phi_stmt_1315_req_0 : boolean;
  signal phi_stmt_1308_ack_0 : boolean;
  signal phi_stmt_1315_ack_0 : boolean;
  signal phi_stmt_1322_ack_0 : boolean;
  signal type_cast_1667_inst_req_0 : boolean;
  signal type_cast_1667_inst_ack_0 : boolean;
  signal type_cast_1667_inst_req_1 : boolean;
  signal type_cast_1667_inst_ack_1 : boolean;
  signal phi_stmt_1662_req_1 : boolean;
  signal type_cast_1659_inst_req_0 : boolean;
  signal type_cast_1659_inst_ack_0 : boolean;
  signal type_cast_1659_inst_req_1 : boolean;
  signal type_cast_1659_inst_ack_1 : boolean;
  signal phi_stmt_1656_req_0 : boolean;
  signal phi_stmt_1649_req_0 : boolean;
  signal type_cast_1665_inst_req_0 : boolean;
  signal type_cast_1665_inst_ack_0 : boolean;
  signal type_cast_1665_inst_req_1 : boolean;
  signal type_cast_1665_inst_ack_1 : boolean;
  signal phi_stmt_1662_req_0 : boolean;
  signal type_cast_1661_inst_req_0 : boolean;
  signal type_cast_1661_inst_ack_0 : boolean;
  signal type_cast_1661_inst_req_1 : boolean;
  signal type_cast_1661_inst_ack_1 : boolean;
  signal phi_stmt_1656_req_1 : boolean;
  signal type_cast_1655_inst_req_0 : boolean;
  signal type_cast_1655_inst_ack_0 : boolean;
  signal type_cast_1655_inst_req_1 : boolean;
  signal type_cast_1655_inst_ack_1 : boolean;
  signal phi_stmt_1649_req_1 : boolean;
  signal phi_stmt_1649_ack_0 : boolean;
  signal phi_stmt_1656_ack_0 : boolean;
  signal phi_stmt_1662_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_B_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_B_CP_3111_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_B_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_B_CP_3111_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_B_CP_3111_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_B_CP_3111_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_B_CP_3111: Block -- control-path 
    signal zeropad3D_B_CP_3111_elements: BooleanArray(134 downto 0);
    -- 
  begin -- 
    zeropad3D_B_CP_3111_elements(0) <= zeropad3D_B_CP_3111_start;
    zeropad3D_B_CP_3111_symbol <= zeropad3D_B_CP_3111_elements(88);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1173/$entry
      -- CP-element group 0: 	 branch_block_stmt_1173/branch_block_stmt_1173__entry__
      -- CP-element group 0: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194__entry__
      -- CP-element group 0: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/$entry
      -- CP-element group 0: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_Sample/rr
      -- 
    rr_3177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(0), ack => RPIPE_Block1_starting_1175_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	134 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1: 	98 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	101 
    -- CP-element group 1: 	102 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_1173/merge_stmt_1648__exit__
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/SplitProtocol/Update/cr
      -- 
    rr_4013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(1), ack => type_cast_1327_inst_req_0); -- 
    cr_4018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(1), ack => type_cast_1327_inst_req_1); -- 
    rr_4036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(1), ack => type_cast_1314_inst_req_0); -- 
    cr_4041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(1), ack => type_cast_1314_inst_req_1); -- 
    rr_4059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(1), ack => type_cast_1318_inst_req_0); -- 
    cr_4064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(1), ack => type_cast_1318_inst_req_1); -- 
    zeropad3D_B_CP_3111_elements(1) <= zeropad3D_B_CP_3111_elements(134);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_Update/cr
      -- 
    ra_3178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1175_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(2)); -- 
    cr_3182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(2), ack => RPIPE_Block1_starting_1175_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1175_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_Sample/rr
      -- 
    ca_3183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1175_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(3)); -- 
    rr_3191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(3), ack => RPIPE_Block1_starting_1178_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_Update/cr
      -- 
    ra_3192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1178_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(4)); -- 
    cr_3196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(4), ack => RPIPE_Block1_starting_1178_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1178_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_Sample/rr
      -- 
    ca_3197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1178_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(5)); -- 
    rr_3205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(5), ack => RPIPE_Block1_starting_1181_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_Update/cr
      -- 
    ra_3206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1181_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(6)); -- 
    cr_3210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(6), ack => RPIPE_Block1_starting_1181_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1181_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_Sample/rr
      -- 
    ca_3211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1181_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(7)); -- 
    rr_3219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(7), ack => RPIPE_Block1_starting_1184_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_Update/cr
      -- 
    ra_3220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1184_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(8)); -- 
    cr_3224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(8), ack => RPIPE_Block1_starting_1184_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1184_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_Sample/rr
      -- 
    ca_3225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1184_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(9)); -- 
    rr_3233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(9), ack => RPIPE_Block1_starting_1187_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_Update/cr
      -- 
    ra_3234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1187_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(10)); -- 
    cr_3238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(10), ack => RPIPE_Block1_starting_1187_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1187_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_Sample/rr
      -- 
    ca_3239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1187_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(11)); -- 
    rr_3247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(11), ack => RPIPE_Block1_starting_1190_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_Update/cr
      -- 
    ra_3248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1190_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(12)); -- 
    cr_3252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(12), ack => RPIPE_Block1_starting_1190_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1190_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_Sample/rr
      -- 
    ca_3253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1190_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(13)); -- 
    rr_3261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(13), ack => RPIPE_Block1_starting_1193_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_Update/cr
      -- 
    ra_3262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1193_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(14)); -- 
    cr_3266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(14), ack => RPIPE_Block1_starting_1193_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	30 
    -- CP-element group 15: 	31 
    -- CP-element group 15:  members (55) 
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194__exit__
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305__entry__
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/$exit
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1176_to_assign_stmt_1194/RPIPE_Block1_starting_1193_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_update_start_
      -- 
    ca_3267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_starting_1193_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(15)); -- 
    cr_3325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1216_inst_req_1); -- 
    cr_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1233_inst_req_1); -- 
    rr_3320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1216_inst_req_0); -- 
    rr_3334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1220_inst_req_0); -- 
    rr_3376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1263_inst_req_0); -- 
    rr_3348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1229_inst_req_0); -- 
    rr_3362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1233_inst_req_0); -- 
    cr_3353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1229_inst_req_1); -- 
    cr_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1263_inst_req_1); -- 
    cr_3339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1220_inst_req_1); -- 
    rr_3278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1198_inst_req_0); -- 
    cr_3283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1198_inst_req_1); -- 
    rr_3292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1208_inst_req_0); -- 
    cr_3297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1208_inst_req_1); -- 
    rr_3306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1212_inst_req_0); -- 
    cr_3311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(15), ack => type_cast_1212_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_Sample/ra
      -- 
    ra_3279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1198_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1198_Update/ca
      -- 
    ca_3284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1198_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_Sample/ra
      -- 
    ra_3293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1208_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	32 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1208_Update/ca
      -- 
    ca_3298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1208_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_Sample/ra
      -- 
    ra_3307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1212_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	32 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1212_Update/ca
      -- 
    ca_3312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1212_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_sample_completed_
      -- 
    ra_3321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1216_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	32 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1216_update_completed_
      -- 
    ca_3326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1216_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_sample_completed_
      -- 
    ra_3335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	32 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1220_Update/ca
      -- 
    ca_3340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_Sample/ra
      -- 
    ra_3349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1229_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	32 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1229_Update/ca
      -- 
    ca_3354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1229_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_Sample/$exit
      -- 
    ra_3363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1233_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1233_update_completed_
      -- 
    ca_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1233_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_Sample/ra
      -- 
    ra_3377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1263_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/type_cast_1263_Update/ca
      -- 
    ca_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1263_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  place  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: 	19 
    -- CP-element group 32: 	21 
    -- CP-element group 32: 	23 
    -- CP-element group 32: 	25 
    -- CP-element group 32: 	27 
    -- CP-element group 32: 	29 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: 	90 
    -- CP-element group 32: 	92 
    -- CP-element group 32: 	93 
    -- CP-element group 32:  members (16) 
      -- CP-element group 32: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305__exit__
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody
      -- CP-element group 32: 	 branch_block_stmt_1173/assign_stmt_1199_to_assign_stmt_1305/$exit
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/$entry
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/$entry
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1308/$entry
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1315/$entry
      -- CP-element group 32: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/$entry
      -- 
    rr_3971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(32), ack => type_cast_1325_inst_req_0); -- 
    cr_3976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(32), ack => type_cast_1325_inst_req_1); -- 
    zeropad3D_B_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(17) & zeropad3D_B_CP_3111_elements(19) & zeropad3D_B_CP_3111_elements(21) & zeropad3D_B_CP_3111_elements(23) & zeropad3D_B_CP_3111_elements(25) & zeropad3D_B_CP_3111_elements(27) & zeropad3D_B_CP_3111_elements(29) & zeropad3D_B_CP_3111_elements(31);
      gj_zeropad3D_B_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	109 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_Sample/$exit
      -- 
    ra_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1332_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(33)); -- 
    -- CP-element group 34:  branch  transition  place  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	109 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (13) 
      -- CP-element group 34: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1173/if_stmt_1359_else_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1173/R_orx_xcond_1360_place
      -- CP-element group 34: 	 branch_block_stmt_1173/if_stmt_1359_dead_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/$exit
      -- CP-element group 34: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1173/if_stmt_1359_eval_test/$entry
      -- CP-element group 34: 	 branch_block_stmt_1173/if_stmt_1359_if_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1173/if_stmt_1359_eval_test/$exit
      -- CP-element group 34: 	 branch_block_stmt_1173/if_stmt_1359_eval_test/branch_req
      -- CP-element group 34: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358__exit__
      -- CP-element group 34: 	 branch_block_stmt_1173/if_stmt_1359__entry__
      -- 
    ca_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1332_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(34)); -- 
    branch_req_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(34), ack => if_stmt_1359_branch_req_0); -- 
    -- CP-element group 35:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (18) 
      -- CP-element group 35: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_1173/if_stmt_1359_if_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_1173/whilex_xbody_lorx_xlhsx_xfalse60
      -- CP-element group 35: 	 branch_block_stmt_1173/if_stmt_1359_if_link/if_choice_transition
      -- CP-element group 35: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/$entry
      -- CP-element group 35: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1173/merge_stmt_1365__exit__
      -- CP-element group 35: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395__entry__
      -- CP-element group 35: 	 branch_block_stmt_1173/whilex_xbody_lorx_xlhsx_xfalse60_PhiReq/$entry
      -- CP-element group 35: 	 branch_block_stmt_1173/whilex_xbody_lorx_xlhsx_xfalse60_PhiReq/$exit
      -- CP-element group 35: 	 branch_block_stmt_1173/merge_stmt_1365_PhiReqMerge
      -- CP-element group 35: 	 branch_block_stmt_1173/merge_stmt_1365_PhiAck/$entry
      -- CP-element group 35: 	 branch_block_stmt_1173/merge_stmt_1365_PhiAck/$exit
      -- CP-element group 35: 	 branch_block_stmt_1173/merge_stmt_1365_PhiAck/dummy
      -- 
    if_choice_transition_3412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1359_branch_ack_1, ack => zeropad3D_B_CP_3111_elements(35)); -- 
    cr_3434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(35), ack => type_cast_1369_inst_req_1); -- 
    rr_3429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(35), ack => type_cast_1369_inst_req_0); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	110 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_1173/if_stmt_1359_else_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_1173/if_stmt_1359_else_link/else_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_1173/whilex_xbody_ifx_xthen
      -- CP-element group 36: 	 branch_block_stmt_1173/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_1173/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_3416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1359_branch_ack_0, ack => zeropad3D_B_CP_3111_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_Sample/$exit
      -- 
    ra_3430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1369_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(37)); -- 
    -- CP-element group 38:  branch  transition  place  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (13) 
      -- CP-element group 38: 	 branch_block_stmt_1173/if_stmt_1396_dead_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_1173/R_orx_xcond190_1397_place
      -- CP-element group 38: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/$exit
      -- CP-element group 38: 	 branch_block_stmt_1173/if_stmt_1396_if_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395/type_cast_1369_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1173/if_stmt_1396_eval_test/$entry
      -- CP-element group 38: 	 branch_block_stmt_1173/if_stmt_1396_eval_test/$exit
      -- CP-element group 38: 	 branch_block_stmt_1173/if_stmt_1396_eval_test/branch_req
      -- CP-element group 38: 	 branch_block_stmt_1173/assign_stmt_1370_to_assign_stmt_1395__exit__
      -- CP-element group 38: 	 branch_block_stmt_1173/if_stmt_1396__entry__
      -- CP-element group 38: 	 branch_block_stmt_1173/if_stmt_1396_else_link/$entry
      -- 
    ca_3435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1369_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(38)); -- 
    branch_req_3443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(38), ack => if_stmt_1396_branch_req_0); -- 
    -- CP-element group 39:  fork  transition  place  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	55 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	58 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	62 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	66 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	70 
    -- CP-element group 39: 	73 
    -- CP-element group 39:  members (46) 
      -- CP-element group 39: 	 branch_block_stmt_1173/if_stmt_1396_if_link/if_choice_transition
      -- CP-element group 39: 	 branch_block_stmt_1173/lorx_xlhsx_xfalse60_ifx_xelse
      -- CP-element group 39: 	 branch_block_stmt_1173/if_stmt_1396_if_link/$exit
      -- CP-element group 39: 	 branch_block_stmt_1173/merge_stmt_1460__exit__
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565__entry__
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_complete/req
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_complete/req
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_1173/lorx_xlhsx_xfalse60_ifx_xelse_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/lorx_xlhsx_xfalse60_ifx_xelse_PhiReq/$exit
      -- CP-element group 39: 	 branch_block_stmt_1173/merge_stmt_1460_PhiReqMerge
      -- CP-element group 39: 	 branch_block_stmt_1173/merge_stmt_1460_PhiAck/$entry
      -- CP-element group 39: 	 branch_block_stmt_1173/merge_stmt_1460_PhiAck/$exit
      -- CP-element group 39: 	 branch_block_stmt_1173/merge_stmt_1460_PhiAck/dummy
      -- 
    if_choice_transition_3448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1396_branch_ack_1, ack => zeropad3D_B_CP_3111_elements(39)); -- 
    rr_3606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(39), ack => type_cast_1464_inst_req_0); -- 
    cr_3611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(39), ack => type_cast_1464_inst_req_1); -- 
    cr_3625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(39), ack => type_cast_1528_inst_req_1); -- 
    req_3656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(39), ack => array_obj_ref_1534_index_offset_req_1); -- 
    req_3671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(39), ack => addr_of_1535_final_reg_req_1); -- 
    cr_3716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(39), ack => ptr_deref_1539_load_0_req_1); -- 
    cr_3735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(39), ack => type_cast_1553_inst_req_1); -- 
    req_3766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(39), ack => array_obj_ref_1559_index_offset_req_1); -- 
    req_3781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(39), ack => addr_of_1560_final_reg_req_1); -- 
    cr_3831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(39), ack => ptr_deref_1563_store_0_req_1); -- 
    -- CP-element group 40:  transition  place  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	110 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1173/lorx_xlhsx_xfalse60_ifx_xthen
      -- CP-element group 40: 	 branch_block_stmt_1173/if_stmt_1396_else_link/else_choice_transition
      -- CP-element group 40: 	 branch_block_stmt_1173/if_stmt_1396_else_link/$exit
      -- CP-element group 40: 	 branch_block_stmt_1173/lorx_xlhsx_xfalse60_ifx_xthen_PhiReq/$entry
      -- CP-element group 40: 	 branch_block_stmt_1173/lorx_xlhsx_xfalse60_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_3452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1396_branch_ack_0, ack => zeropad3D_B_CP_3111_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	110 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_sample_completed_
      -- 
    ra_3466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	110 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_Update/$exit
      -- 
    ca_3471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	110 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_Sample/ra
      -- 
    ra_3480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	110 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_Update/ca
      -- 
    ca_3485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_Sample/rr
      -- CP-element group 45: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_sample_start_
      -- 
    rr_3493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(45), ack => type_cast_1445_inst_req_0); -- 
    zeropad3D_B_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(42) & zeropad3D_B_CP_3111_elements(44);
      gj_zeropad3D_B_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_Sample/$exit
      -- 
    ra_3494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1445_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	110 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (16) 
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_scale_1/scale_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_scale_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_scale_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_resize_1/index_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_scale_1/scale_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_resized_1
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_scaled_1
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_computed_1
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_resize_1/index_resize_req
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_resize_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_index_resize_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_final_index_sum_regn_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_final_index_sum_regn_Sample/req
      -- 
    ca_3499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1445_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(47)); -- 
    req_3524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(47), ack => array_obj_ref_1451_index_offset_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	54 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_final_index_sum_regn_sample_complete
      -- CP-element group 48: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_final_index_sum_regn_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_final_index_sum_regn_Sample/ack
      -- 
    ack_3525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1451_index_offset_ack_0, ack => zeropad3D_B_CP_3111_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	110 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (11) 
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_offset_calculated
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_final_index_sum_regn_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_final_index_sum_regn_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_request/$entry
      -- CP-element group 49: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_request/req
      -- 
    ack_3530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1451_index_offset_ack_1, ack => zeropad3D_B_CP_3111_elements(49)); -- 
    req_3539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(49), ack => addr_of_1452_final_reg_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_request/$exit
      -- CP-element group 50: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_request/ack
      -- 
    ack_3540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1452_final_reg_ack_0, ack => zeropad3D_B_CP_3111_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	110 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (28) 
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_complete/ack
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_base_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_word_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_base_address_resized
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_base_addr_resize/$entry
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_base_addr_resize/$exit
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_base_addr_resize/base_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_base_addr_resize/base_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_word_addrgen/$entry
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_word_addrgen/$exit
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_word_addrgen/root_register_req
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_word_addrgen/root_register_ack
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/ptr_deref_1455_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/ptr_deref_1455_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/ptr_deref_1455_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/ptr_deref_1455_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/word_access_start/word_0/rr
      -- 
    ack_3545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1452_final_reg_ack_1, ack => zeropad3D_B_CP_3111_elements(51)); -- 
    rr_3583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(51), ack => ptr_deref_1455_store_0_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Sample/word_access_start/word_0/ra
      -- 
    ra_3584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1455_store_0_ack_0, ack => zeropad3D_B_CP_3111_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	110 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Update/word_access_complete/word_0/ca
      -- 
    ca_3595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1455_store_0_ack_1, ack => zeropad3D_B_CP_3111_elements(53)); -- 
    -- CP-element group 54:  join  transition  place  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	48 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	111 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/$exit
      -- CP-element group 54: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458__exit__
      -- CP-element group 54: 	 branch_block_stmt_1173/ifx_xthen_ifx_xend
      -- CP-element group 54: 	 branch_block_stmt_1173/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_1173/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(48) & zeropad3D_B_CP_3111_elements(53);
      gj_zeropad3D_B_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	39 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_Sample/ra
      -- 
    ra_3607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1464_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	65 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1464_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_Sample/rr
      -- 
    ca_3612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1464_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(56)); -- 
    rr_3620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(56), ack => type_cast_1528_inst_req_0); -- 
    rr_3730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(56), ack => type_cast_1553_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_Sample/ra
      -- 
    ra_3621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1528_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	39 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (16) 
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1528_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_final_index_sum_regn_Sample/req
      -- 
    ca_3626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1528_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(58)); -- 
    req_3651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(58), ack => array_obj_ref_1534_index_offset_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	74 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_final_index_sum_regn_Sample/ack
      -- 
    ack_3652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1534_index_offset_ack_0, ack => zeropad3D_B_CP_3111_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1534_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_request/req
      -- 
    ack_3657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1534_index_offset_ack_1, ack => zeropad3D_B_CP_3111_elements(60)); -- 
    req_3666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(60), ack => addr_of_1535_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_request/ack
      -- 
    ack_3667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1535_final_reg_ack_0, ack => zeropad3D_B_CP_3111_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	39 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (24) 
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1535_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Sample/word_access_start/word_0/rr
      -- 
    ack_3672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1535_final_reg_ack_1, ack => zeropad3D_B_CP_3111_elements(62)); -- 
    rr_3705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(62), ack => ptr_deref_1539_load_0_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Sample/word_access_start/word_0/ra
      -- 
    ra_3706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1539_load_0_ack_0, ack => zeropad3D_B_CP_3111_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	71 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/ptr_deref_1539_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/ptr_deref_1539_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/ptr_deref_1539_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1539_Update/ptr_deref_1539_Merge/merge_ack
      -- 
    ca_3717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1539_load_0_ack_1, ack => zeropad3D_B_CP_3111_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	56 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_Sample/ra
      -- 
    ra_3731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1553_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	39 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/type_cast_1553_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_resized_1
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_scaled_1
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_computed_1
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_resize_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_resize_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_resize_1/index_resize_req
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_resize_1/index_resize_ack
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_scale_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_scale_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_scale_1/scale_rename_req
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_index_scale_1/scale_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_final_index_sum_regn_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_final_index_sum_regn_Sample/req
      -- 
    ca_3736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1553_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(66)); -- 
    req_3761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(66), ack => array_obj_ref_1559_index_offset_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	74 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_final_index_sum_regn_sample_complete
      -- CP-element group 67: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_final_index_sum_regn_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_final_index_sum_regn_Sample/ack
      -- 
    ack_3762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1559_index_offset_ack_0, ack => zeropad3D_B_CP_3111_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (11) 
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_offset_calculated
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_final_index_sum_regn_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_final_index_sum_regn_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/array_obj_ref_1559_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_request/$entry
      -- CP-element group 68: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_request/req
      -- 
    ack_3767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1559_index_offset_ack_1, ack => zeropad3D_B_CP_3111_elements(68)); -- 
    req_3776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(68), ack => addr_of_1560_final_reg_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_request/$exit
      -- CP-element group 69: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_request/ack
      -- 
    ack_3777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1560_final_reg_ack_0, ack => zeropad3D_B_CP_3111_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	39 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (19) 
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/addr_of_1560_complete/ack
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_base_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_word_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_base_address_resized
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_base_addr_resize/$entry
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_base_addr_resize/$exit
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_base_addr_resize/base_resize_req
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_base_addr_resize/base_resize_ack
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_word_addrgen/$entry
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_word_addrgen/$exit
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_word_addrgen/root_register_req
      -- CP-element group 70: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_word_addrgen/root_register_ack
      -- 
    ack_3782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1560_final_reg_ack_1, ack => zeropad3D_B_CP_3111_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	64 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/ptr_deref_1563_Split/$entry
      -- CP-element group 71: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/ptr_deref_1563_Split/$exit
      -- CP-element group 71: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/ptr_deref_1563_Split/split_req
      -- CP-element group 71: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/ptr_deref_1563_Split/split_ack
      -- CP-element group 71: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/word_access_start/$entry
      -- CP-element group 71: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/word_access_start/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/word_access_start/word_0/rr
      -- 
    rr_3820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(71), ack => ptr_deref_1563_store_0_req_0); -- 
    zeropad3D_B_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(64) & zeropad3D_B_CP_3111_elements(70);
      gj_zeropad3D_B_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/word_access_start/$exit
      -- CP-element group 72: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/word_access_start/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Sample/word_access_start/word_0/ra
      -- 
    ra_3821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1563_store_0_ack_0, ack => zeropad3D_B_CP_3111_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	39 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Update/word_access_complete/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/ptr_deref_1563_Update/word_access_complete/word_0/ca
      -- 
    ca_3832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1563_store_0_ack_1, ack => zeropad3D_B_CP_3111_elements(73)); -- 
    -- CP-element group 74:  join  transition  place  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	59 
    -- CP-element group 74: 	67 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	111 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565__exit__
      -- CP-element group 74: 	 branch_block_stmt_1173/ifx_xelse_ifx_xend
      -- CP-element group 74: 	 branch_block_stmt_1173/assign_stmt_1465_to_assign_stmt_1565/$exit
      -- CP-element group 74: 	 branch_block_stmt_1173/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_1173/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(59) & zeropad3D_B_CP_3111_elements(67) & zeropad3D_B_CP_3111_elements(73);
      gj_zeropad3D_B_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	111 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_Sample/ra
      -- 
    ra_3844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1571_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(75)); -- 
    -- CP-element group 76:  branch  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	111 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (13) 
      -- CP-element group 76: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585__exit__
      -- CP-element group 76: 	 branch_block_stmt_1173/if_stmt_1586__entry__
      -- CP-element group 76: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/$exit
      -- CP-element group 76: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_1173/if_stmt_1586_dead_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_1173/if_stmt_1586_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_1173/if_stmt_1586_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_1173/if_stmt_1586_eval_test/branch_req
      -- CP-element group 76: 	 branch_block_stmt_1173/R_cmp144_1587_place
      -- CP-element group 76: 	 branch_block_stmt_1173/if_stmt_1586_if_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_1173/if_stmt_1586_else_link/$entry
      -- 
    ca_3849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1571_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(76)); -- 
    branch_req_3857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(76), ack => if_stmt_1586_branch_req_0); -- 
    -- CP-element group 77:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	120 
    -- CP-element group 77: 	121 
    -- CP-element group 77: 	123 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	126 
    -- CP-element group 77: 	127 
    -- CP-element group 77:  members (40) 
      -- CP-element group 77: 	 branch_block_stmt_1173/merge_stmt_1592__exit__
      -- CP-element group 77: 	 branch_block_stmt_1173/assign_stmt_1598__entry__
      -- CP-element group 77: 	 branch_block_stmt_1173/assign_stmt_1598__exit__
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184
      -- CP-element group 77: 	 branch_block_stmt_1173/if_stmt_1586_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_1173/if_stmt_1586_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xend_ifx_xthen146
      -- CP-element group 77: 	 branch_block_stmt_1173/assign_stmt_1598/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/assign_stmt_1598/$exit
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xend_ifx_xthen146_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xend_ifx_xthen146_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_1173/merge_stmt_1592_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_1173/merge_stmt_1592_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/merge_stmt_1592_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_1173/merge_stmt_1592_PhiAck/dummy
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1586_branch_ack_1, ack => zeropad3D_B_CP_3111_elements(77)); -- 
    rr_4219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(77), ack => type_cast_1665_inst_req_0); -- 
    cr_4224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(77), ack => type_cast_1665_inst_req_1); -- 
    rr_4242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(77), ack => type_cast_1661_inst_req_0); -- 
    cr_4247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(77), ack => type_cast_1661_inst_req_1); -- 
    rr_4265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(77), ack => type_cast_1655_inst_req_0); -- 
    cr_4270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(77), ack => type_cast_1655_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	84 
    -- CP-element group 78:  members (24) 
      -- CP-element group 78: 	 branch_block_stmt_1173/merge_stmt_1600__exit__
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641__entry__
      -- CP-element group 78: 	 branch_block_stmt_1173/if_stmt_1586_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_1173/if_stmt_1586_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_1173/ifx_xend_ifx_xelse151
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/$entry
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_1173/ifx_xend_ifx_xelse151_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1173/ifx_xend_ifx_xelse151_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1173/merge_stmt_1600_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1173/merge_stmt_1600_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1173/merge_stmt_1600_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1173/merge_stmt_1600_PhiAck/dummy
      -- 
    else_choice_transition_3866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1586_branch_ack_0, ack => zeropad3D_B_CP_3111_elements(78)); -- 
    rr_3882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(78), ack => type_cast_1610_inst_req_0); -- 
    cr_3887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(78), ack => type_cast_1610_inst_req_1); -- 
    cr_3901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(78), ack => type_cast_1619_inst_req_1); -- 
    cr_3915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(78), ack => type_cast_1635_inst_req_1); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_Sample/ra
      -- 
    ra_3883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1610_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1610_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_Sample/rr
      -- 
    ca_3888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1610_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(80)); -- 
    rr_3896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(80), ack => type_cast_1619_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_Sample/ra
      -- 
    ra_3897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1619_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1619_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_Sample/rr
      -- 
    ca_3902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1619_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(82)); -- 
    rr_3910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(82), ack => type_cast_1635_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_Sample/ra
      -- 
    ra_3911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1635_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(83)); -- 
    -- CP-element group 84:  branch  transition  place  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	78 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (13) 
      -- CP-element group 84: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641__exit__
      -- CP-element group 84: 	 branch_block_stmt_1173/if_stmt_1642__entry__
      -- CP-element group 84: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/$exit
      -- CP-element group 84: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_1173/assign_stmt_1606_to_assign_stmt_1641/type_cast_1635_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_1173/if_stmt_1642_dead_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_1173/if_stmt_1642_eval_test/$entry
      -- CP-element group 84: 	 branch_block_stmt_1173/if_stmt_1642_eval_test/$exit
      -- CP-element group 84: 	 branch_block_stmt_1173/if_stmt_1642_eval_test/branch_req
      -- CP-element group 84: 	 branch_block_stmt_1173/R_cmp176_1643_place
      -- CP-element group 84: 	 branch_block_stmt_1173/if_stmt_1642_if_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_1173/if_stmt_1642_else_link/$entry
      -- 
    ca_3916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1635_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(84)); -- 
    branch_req_3924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(84), ack => if_stmt_1642_branch_req_0); -- 
    -- CP-element group 85:  transition  place  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (15) 
      -- CP-element group 85: 	 branch_block_stmt_1173/merge_stmt_1670__exit__
      -- CP-element group 85: 	 branch_block_stmt_1173/assign_stmt_1675__entry__
      -- CP-element group 85: 	 branch_block_stmt_1173/if_stmt_1642_if_link/$exit
      -- CP-element group 85: 	 branch_block_stmt_1173/if_stmt_1642_if_link/if_choice_transition
      -- CP-element group 85: 	 branch_block_stmt_1173/ifx_xelse151_whilex_xend
      -- CP-element group 85: 	 branch_block_stmt_1173/assign_stmt_1675/$entry
      -- CP-element group 85: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_1173/ifx_xelse151_whilex_xend_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_1173/ifx_xelse151_whilex_xend_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1173/merge_stmt_1670_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_1173/merge_stmt_1670_PhiAck/$entry
      -- CP-element group 85: 	 branch_block_stmt_1173/merge_stmt_1670_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_1173/merge_stmt_1670_PhiAck/dummy
      -- 
    if_choice_transition_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1642_branch_ack_1, ack => zeropad3D_B_CP_3111_elements(85)); -- 
    req_3946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(85), ack => WPIPE_Block1_complete_1672_inst_req_0); -- 
    -- CP-element group 86:  fork  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	112 
    -- CP-element group 86: 	113 
    -- CP-element group 86: 	115 
    -- CP-element group 86: 	116 
    -- CP-element group 86: 	118 
    -- CP-element group 86:  members (22) 
      -- CP-element group 86: 	 branch_block_stmt_1173/if_stmt_1642_else_link/$exit
      -- CP-element group 86: 	 branch_block_stmt_1173/if_stmt_1642_else_link/else_choice_transition
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1649/$entry
      -- CP-element group 86: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/$entry
      -- 
    else_choice_transition_3933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1642_branch_ack_0, ack => zeropad3D_B_CP_3111_elements(86)); -- 
    rr_4162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(86), ack => type_cast_1667_inst_req_0); -- 
    cr_4167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(86), ack => type_cast_1667_inst_req_1); -- 
    rr_4185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(86), ack => type_cast_1659_inst_req_0); -- 
    cr_4190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(86), ack => type_cast_1659_inst_req_1); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_Update/req
      -- 
    ack_3947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_complete_1672_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(87)); -- 
    req_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(87), ack => WPIPE_Block1_complete_1672_inst_req_1); -- 
    -- CP-element group 88:  transition  place  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 $exit
      -- CP-element group 88: 	 branch_block_stmt_1173/$exit
      -- CP-element group 88: 	 branch_block_stmt_1173/branch_block_stmt_1173__exit__
      -- CP-element group 88: 	 branch_block_stmt_1173/assign_stmt_1675__exit__
      -- CP-element group 88: 	 branch_block_stmt_1173/return__
      -- CP-element group 88: 	 branch_block_stmt_1173/merge_stmt_1677__exit__
      -- CP-element group 88: 	 branch_block_stmt_1173/assign_stmt_1675/$exit
      -- CP-element group 88: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1173/assign_stmt_1675/WPIPE_Block1_complete_1672_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_1173/return___PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_1173/return___PhiReq/$exit
      -- CP-element group 88: 	 branch_block_stmt_1173/merge_stmt_1677_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_1173/merge_stmt_1677_PhiAck/$entry
      -- CP-element group 88: 	 branch_block_stmt_1173/merge_stmt_1677_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_1173/merge_stmt_1677_PhiAck/dummy
      -- 
    ack_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_complete_1672_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/SplitProtocol/Sample/ra
      -- 
    ra_3972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	32 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/SplitProtocol/Update/ca
      -- 
    ca_3977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/$exit
      -- CP-element group 91: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/$exit
      -- CP-element group 91: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1325/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_req
      -- 
    phi_stmt_1322_req_3978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1322_req_3978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(91), ack => phi_stmt_1322_req_0); -- 
    zeropad3D_B_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(89) & zeropad3D_B_CP_3111_elements(90);
      gj_zeropad3D_B_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  output  delay-element  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	32 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1308/$exit
      -- CP-element group 92: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1312_konst_delay_trans
      -- CP-element group 92: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_req
      -- 
    phi_stmt_1308_req_3986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1308_req_3986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(92), ack => phi_stmt_1308_req_0); -- 
    -- Element group zeropad3D_B_CP_3111_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => zeropad3D_B_CP_3111_elements(32), ack => zeropad3D_B_CP_3111_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  transition  output  delay-element  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	32 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1315/$exit
      -- CP-element group 93: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1321_konst_delay_trans
      -- CP-element group 93: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_req
      -- 
    phi_stmt_1315_req_3994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1315_req_3994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(93), ack => phi_stmt_1315_req_1); -- 
    -- Element group zeropad3D_B_CP_3111_elements(93) is a control-delay.
    cp_element_93_delay: control_delay_element  generic map(name => " 93_delay", delay_value => 1)  port map(req => zeropad3D_B_CP_3111_elements(32), ack => zeropad3D_B_CP_3111_elements(93), clk => clk, reset =>reset);
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	105 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_1173/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(91) & zeropad3D_B_CP_3111_elements(92) & zeropad3D_B_CP_3111_elements(93);
      gj_zeropad3D_B_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/SplitProtocol/Sample/ra
      -- 
    ra_4014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1327_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/SplitProtocol/Update/ca
      -- 
    ca_4019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1327_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	104 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/$exit
      -- CP-element group 97: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/$exit
      -- CP-element group 97: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_sources/type_cast_1327/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1322/phi_stmt_1322_req
      -- 
    phi_stmt_1322_req_4020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1322_req_4020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(97), ack => phi_stmt_1322_req_1); -- 
    zeropad3D_B_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_B_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(95) & zeropad3D_B_CP_3111_elements(96);
      gj_zeropad3D_B_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	1 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/SplitProtocol/Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/SplitProtocol/Sample/ra
      -- 
    ra_4037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1314_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/SplitProtocol/Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/SplitProtocol/Update/ca
      -- 
    ca_4042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1314_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/$exit
      -- CP-element group 100: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/$exit
      -- CP-element group 100: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_sources/type_cast_1314/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1308/phi_stmt_1308_req
      -- 
    phi_stmt_1308_req_4043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1308_req_4043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(100), ack => phi_stmt_1308_req_1); -- 
    zeropad3D_B_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(98) & zeropad3D_B_CP_3111_elements(99);
      gj_zeropad3D_B_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	1 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/SplitProtocol/Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/SplitProtocol/Sample/ra
      -- 
    ra_4060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1318_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/SplitProtocol/Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/SplitProtocol/Update/ca
      -- 
    ca_4065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1318_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/$exit
      -- CP-element group 103: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/$exit
      -- CP-element group 103: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/type_cast_1318/SplitProtocol/$exit
      -- CP-element group 103: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_1315/phi_stmt_1315_req
      -- 
    phi_stmt_1315_req_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1315_req_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(103), ack => phi_stmt_1315_req_0); -- 
    zeropad3D_B_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(101) & zeropad3D_B_CP_3111_elements(102);
      gj_zeropad3D_B_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	97 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1173/ifx_xend184_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(97) & zeropad3D_B_CP_3111_elements(100) & zeropad3D_B_CP_3111_elements(103);
      gj_zeropad3D_B_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  merge  fork  transition  place  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	94 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1173/merge_stmt_1307_PhiReqMerge
      -- CP-element group 105: 	 branch_block_stmt_1173/merge_stmt_1307_PhiAck/$entry
      -- 
    zeropad3D_B_CP_3111_elements(105) <= OrReduce(zeropad3D_B_CP_3111_elements(94) & zeropad3D_B_CP_3111_elements(104));
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	109 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1173/merge_stmt_1307_PhiAck/phi_stmt_1308_ack
      -- 
    phi_stmt_1308_ack_4071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1308_ack_0, ack => zeropad3D_B_CP_3111_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_1173/merge_stmt_1307_PhiAck/phi_stmt_1315_ack
      -- 
    phi_stmt_1315_ack_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1315_ack_0, ack => zeropad3D_B_CP_3111_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1173/merge_stmt_1307_PhiAck/phi_stmt_1322_ack
      -- 
    phi_stmt_1322_ack_4073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1322_ack_0, ack => zeropad3D_B_CP_3111_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  place  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	106 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	34 
    -- CP-element group 109: 	33 
    -- CP-element group 109:  members (10) 
      -- CP-element group 109: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/type_cast_1332_Update/cr
      -- CP-element group 109: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358/$entry
      -- CP-element group 109: 	 branch_block_stmt_1173/merge_stmt_1307__exit__
      -- CP-element group 109: 	 branch_block_stmt_1173/assign_stmt_1333_to_assign_stmt_1358__entry__
      -- CP-element group 109: 	 branch_block_stmt_1173/merge_stmt_1307_PhiAck/$exit
      -- 
    rr_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(109), ack => type_cast_1332_inst_req_0); -- 
    cr_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(109), ack => type_cast_1332_inst_req_1); -- 
    zeropad3D_B_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(106) & zeropad3D_B_CP_3111_elements(107) & zeropad3D_B_CP_3111_elements(108);
      gj_zeropad3D_B_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  merge  fork  transition  place  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	40 
    -- CP-element group 110: 	36 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	42 
    -- CP-element group 110: 	49 
    -- CP-element group 110: 	51 
    -- CP-element group 110: 	47 
    -- CP-element group 110: 	44 
    -- CP-element group 110: 	53 
    -- CP-element group 110: 	43 
    -- CP-element group 110: 	41 
    -- CP-element group 110:  members (33) 
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_final_index_sum_regn_update_start
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1445_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1406_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/type_cast_1411_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_final_index_sum_regn_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/array_obj_ref_1451_final_index_sum_regn_Update/req
      -- CP-element group 110: 	 branch_block_stmt_1173/merge_stmt_1402__exit__
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458__entry__
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/addr_of_1452_complete/req
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Update/word_access_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Update/word_access_complete/word_0/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/assign_stmt_1407_to_assign_stmt_1458/ptr_deref_1455_Update/word_access_complete/word_0/cr
      -- CP-element group 110: 	 branch_block_stmt_1173/merge_stmt_1402_PhiReqMerge
      -- CP-element group 110: 	 branch_block_stmt_1173/merge_stmt_1402_PhiAck/$entry
      -- CP-element group 110: 	 branch_block_stmt_1173/merge_stmt_1402_PhiAck/$exit
      -- CP-element group 110: 	 branch_block_stmt_1173/merge_stmt_1402_PhiAck/dummy
      -- 
    rr_3465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(110), ack => type_cast_1406_inst_req_0); -- 
    cr_3498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(110), ack => type_cast_1445_inst_req_1); -- 
    rr_3479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(110), ack => type_cast_1411_inst_req_0); -- 
    cr_3484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(110), ack => type_cast_1411_inst_req_1); -- 
    cr_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(110), ack => type_cast_1406_inst_req_1); -- 
    req_3529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(110), ack => array_obj_ref_1451_index_offset_req_1); -- 
    req_3544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(110), ack => addr_of_1452_final_reg_req_1); -- 
    cr_3594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(110), ack => ptr_deref_1455_store_0_req_1); -- 
    zeropad3D_B_CP_3111_elements(110) <= OrReduce(zeropad3D_B_CP_3111_elements(40) & zeropad3D_B_CP_3111_elements(36));
    -- CP-element group 111:  merge  fork  transition  place  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	54 
    -- CP-element group 111: 	74 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	75 
    -- CP-element group 111: 	76 
    -- CP-element group 111:  members (13) 
      -- CP-element group 111: 	 branch_block_stmt_1173/merge_stmt_1567__exit__
      -- CP-element group 111: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585__entry__
      -- CP-element group 111: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/$entry
      -- CP-element group 111: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1173/assign_stmt_1572_to_assign_stmt_1585/type_cast_1571_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_1173/merge_stmt_1567_PhiReqMerge
      -- CP-element group 111: 	 branch_block_stmt_1173/merge_stmt_1567_PhiAck/$entry
      -- CP-element group 111: 	 branch_block_stmt_1173/merge_stmt_1567_PhiAck/$exit
      -- CP-element group 111: 	 branch_block_stmt_1173/merge_stmt_1567_PhiAck/dummy
      -- 
    rr_3843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(111), ack => type_cast_1571_inst_req_0); -- 
    cr_3848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(111), ack => type_cast_1571_inst_req_1); -- 
    zeropad3D_B_CP_3111_elements(111) <= OrReduce(zeropad3D_B_CP_3111_elements(54) & zeropad3D_B_CP_3111_elements(74));
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	86 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/SplitProtocol/Sample/ra
      -- 
    ra_4163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1667_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	86 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/SplitProtocol/Update/ca
      -- 
    ca_4168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1667_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	119 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/$exit
      -- CP-element group 114: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/$exit
      -- CP-element group 114: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1667/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_req
      -- 
    phi_stmt_1662_req_4169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1662_req_4169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(114), ack => phi_stmt_1662_req_1); -- 
    zeropad3D_B_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(112) & zeropad3D_B_CP_3111_elements(113);
      gj_zeropad3D_B_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	86 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/SplitProtocol/Sample/ra
      -- 
    ra_4186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1659_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	86 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/SplitProtocol/Update/ca
      -- 
    ca_4191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1659_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/$exit
      -- CP-element group 117: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/$exit
      -- CP-element group 117: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1659/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_req
      -- 
    phi_stmt_1656_req_4192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1656_req_4192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(117), ack => phi_stmt_1656_req_0); -- 
    zeropad3D_B_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(115) & zeropad3D_B_CP_3111_elements(116);
      gj_zeropad3D_B_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  output  delay-element  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	86 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1649/$exit
      -- CP-element group 118: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1653_konst_delay_trans
      -- CP-element group 118: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_req
      -- 
    phi_stmt_1649_req_4200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1649_req_4200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(118), ack => phi_stmt_1649_req_0); -- 
    -- Element group zeropad3D_B_CP_3111_elements(118) is a control-delay.
    cp_element_118_delay: control_delay_element  generic map(name => " 118_delay", delay_value => 1)  port map(req => zeropad3D_B_CP_3111_elements(86), ack => zeropad3D_B_CP_3111_elements(118), clk => clk, reset =>reset);
    -- CP-element group 119:  join  transition  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	114 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	130 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1173/ifx_xelse151_ifx_xend184_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(114) & zeropad3D_B_CP_3111_elements(117) & zeropad3D_B_CP_3111_elements(118);
      gj_zeropad3D_B_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	77 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/SplitProtocol/Sample/ra
      -- 
    ra_4220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1665_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	77 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/SplitProtocol/Update/ca
      -- 
    ca_4225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1665_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	129 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/$exit
      -- CP-element group 122: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/$exit
      -- CP-element group 122: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_sources/type_cast_1665/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1662/phi_stmt_1662_req
      -- 
    phi_stmt_1662_req_4226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1662_req_4226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(122), ack => phi_stmt_1662_req_0); -- 
    zeropad3D_B_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(120) & zeropad3D_B_CP_3111_elements(121);
      gj_zeropad3D_B_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	77 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/SplitProtocol/Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/SplitProtocol/Sample/ra
      -- 
    ra_4243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1661_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/SplitProtocol/Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/SplitProtocol/Update/ca
      -- 
    ca_4248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1661_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	129 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/$exit
      -- CP-element group 125: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/$exit
      -- CP-element group 125: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/$exit
      -- CP-element group 125: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_sources/type_cast_1661/SplitProtocol/$exit
      -- CP-element group 125: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1656/phi_stmt_1656_req
      -- 
    phi_stmt_1656_req_4249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1656_req_4249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(125), ack => phi_stmt_1656_req_1); -- 
    zeropad3D_B_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(123) & zeropad3D_B_CP_3111_elements(124);
      gj_zeropad3D_B_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	77 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/SplitProtocol/Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/SplitProtocol/Sample/ra
      -- 
    ra_4266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1655_inst_ack_0, ack => zeropad3D_B_CP_3111_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	77 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/SplitProtocol/Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/SplitProtocol/Update/ca
      -- 
    ca_4271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1655_inst_ack_1, ack => zeropad3D_B_CP_3111_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/$exit
      -- CP-element group 128: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/$exit
      -- CP-element group 128: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/$exit
      -- CP-element group 128: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_sources/type_cast_1655/SplitProtocol/$exit
      -- CP-element group 128: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/phi_stmt_1649/phi_stmt_1649_req
      -- 
    phi_stmt_1649_req_4272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1649_req_4272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_B_CP_3111_elements(128), ack => phi_stmt_1649_req_1); -- 
    zeropad3D_B_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(126) & zeropad3D_B_CP_3111_elements(127);
      gj_zeropad3D_B_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	122 
    -- CP-element group 129: 	125 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1173/ifx_xthen146_ifx_xend184_PhiReq/$exit
      -- 
    zeropad3D_B_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(122) & zeropad3D_B_CP_3111_elements(125) & zeropad3D_B_CP_3111_elements(128);
      gj_zeropad3D_B_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  fork  transition  place  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	119 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	132 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_1173/merge_stmt_1648_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_1173/merge_stmt_1648_PhiAck/$entry
      -- 
    zeropad3D_B_CP_3111_elements(130) <= OrReduce(zeropad3D_B_CP_3111_elements(119) & zeropad3D_B_CP_3111_elements(129));
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	134 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1173/merge_stmt_1648_PhiAck/phi_stmt_1649_ack
      -- 
    phi_stmt_1649_ack_4277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1649_ack_0, ack => zeropad3D_B_CP_3111_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_1173/merge_stmt_1648_PhiAck/phi_stmt_1656_ack
      -- 
    phi_stmt_1656_ack_4278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1656_ack_0, ack => zeropad3D_B_CP_3111_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_1173/merge_stmt_1648_PhiAck/phi_stmt_1662_ack
      -- 
    phi_stmt_1662_ack_4279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1662_ack_0, ack => zeropad3D_B_CP_3111_elements(133)); -- 
    -- CP-element group 134:  join  transition  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	131 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	1 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_1173/merge_stmt_1648_PhiAck/$exit
      -- 
    zeropad3D_B_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_B_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_B_CP_3111_elements(131) & zeropad3D_B_CP_3111_elements(132) & zeropad3D_B_CP_3111_elements(133);
      gj_zeropad3D_B_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_B_CP_3111_elements(134), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1247_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1303_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1439_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1522_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1547_wire : std_logic_vector(31 downto 0);
    signal R_idxprom131_1533_resized : std_logic_vector(13 downto 0);
    signal R_idxprom131_1533_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom136_1558_resized : std_logic_vector(13 downto 0);
    signal R_idxprom136_1558_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1450_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1450_scaled : std_logic_vector(13 downto 0);
    signal add103_1490 : std_logic_vector(31 downto 0);
    signal add112_1495 : std_logic_vector(31 downto 0);
    signal add122_1510 : std_logic_vector(31 downto 0);
    signal add128_1515 : std_logic_vector(31 downto 0);
    signal add141_1578 : std_logic_vector(31 downto 0);
    signal add149_1598 : std_logic_vector(15 downto 0);
    signal add159_1260 : std_logic_vector(31 downto 0);
    signal add175_1275 : std_logic_vector(31 downto 0);
    signal add74_1285 : std_logic_vector(31 downto 0);
    signal add85_1427 : std_logic_vector(31 downto 0);
    signal add91_1432 : std_logic_vector(31 downto 0);
    signal add_1280 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1451_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1451_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1451_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1451_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1451_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1451_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1534_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1534_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1534_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1534_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1534_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1534_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1559_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1559_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1559_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1559_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1559_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1559_root_address : std_logic_vector(13 downto 0);
    signal arrayidx132_1536 : std_logic_vector(31 downto 0);
    signal arrayidx137_1561 : std_logic_vector(31 downto 0);
    signal arrayidx_1453 : std_logic_vector(31 downto 0);
    signal call1_1179 : std_logic_vector(7 downto 0);
    signal call2_1182 : std_logic_vector(7 downto 0);
    signal call3_1185 : std_logic_vector(7 downto 0);
    signal call4_1188 : std_logic_vector(7 downto 0);
    signal call5_1191 : std_logic_vector(7 downto 0);
    signal call6_1194 : std_logic_vector(7 downto 0);
    signal call_1176 : std_logic_vector(7 downto 0);
    signal cmp144_1585 : std_logic_vector(0 downto 0);
    signal cmp160_1616 : std_logic_vector(0 downto 0);
    signal cmp176_1641 : std_logic_vector(0 downto 0);
    signal cmp58_1353 : std_logic_vector(0 downto 0);
    signal cmp65_1377 : std_logic_vector(0 downto 0);
    signal cmp65x_xnot_1383 : std_logic_vector(0 downto 0);
    signal cmp75_1390 : std_logic_vector(0 downto 0);
    signal cmp_1340 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_1346 : std_logic_vector(0 downto 0);
    signal conv105_1305 : std_logic_vector(31 downto 0);
    signal conv140_1572 : std_logic_vector(31 downto 0);
    signal conv154_1611 : std_logic_vector(31 downto 0);
    signal conv168_1636 : std_logic_vector(31 downto 0);
    signal conv170_1264 : std_logic_vector(31 downto 0);
    signal conv32_1209 : std_logic_vector(31 downto 0);
    signal conv34_1213 : std_logic_vector(31 downto 0);
    signal conv38_1217 : std_logic_vector(31 downto 0);
    signal conv40_1221 : std_logic_vector(31 downto 0);
    signal conv47_1333 : std_logic_vector(31 downto 0);
    signal conv49_1230 : std_logic_vector(31 downto 0);
    signal conv62_1370 : std_logic_vector(31 downto 0);
    signal conv79_1407 : std_logic_vector(31 downto 0);
    signal conv81_1234 : std_logic_vector(31 downto 0);
    signal conv83_1412 : std_logic_vector(31 downto 0);
    signal conv87_1249 : std_logic_vector(31 downto 0);
    signal conv95_1465 : std_logic_vector(31 downto 0);
    signal conv_1199 : std_logic_vector(15 downto 0);
    signal div171_1270 : std_logic_vector(31 downto 0);
    signal div_1205 : std_logic_vector(15 downto 0);
    signal idxprom131_1529 : std_logic_vector(63 downto 0);
    signal idxprom136_1554 : std_logic_vector(63 downto 0);
    signal idxprom_1446 : std_logic_vector(63 downto 0);
    signal inc165_1620 : std_logic_vector(15 downto 0);
    signal inc165x_xix_x2_1625 : std_logic_vector(15 downto 0);
    signal inc_1606 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_1656 : std_logic_vector(15 downto 0);
    signal ix_x2_1315 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_1662 : std_logic_vector(15 downto 0);
    signal jx_x1_1322 : std_logic_vector(15 downto 0);
    signal jx_x2_1631 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_1649 : std_logic_vector(15 downto 0);
    signal kx_x1_1308 : std_logic_vector(15 downto 0);
    signal mul102_1475 : std_logic_vector(31 downto 0);
    signal mul111_1485 : std_logic_vector(31 downto 0);
    signal mul121_1500 : std_logic_vector(31 downto 0);
    signal mul127_1505 : std_logic_vector(31 downto 0);
    signal mul41_1226 : std_logic_vector(31 downto 0);
    signal mul84_1417 : std_logic_vector(31 downto 0);
    signal mul90_1422 : std_logic_vector(31 downto 0);
    signal mul_1291 : std_logic_vector(31 downto 0);
    signal orx_xcond190_1395 : std_logic_vector(0 downto 0);
    signal orx_xcond_1358 : std_logic_vector(0 downto 0);
    signal ptr_deref_1455_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1455_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1455_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1455_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1455_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1455_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1539_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1539_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1539_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1539_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1539_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1563_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1563_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1563_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1563_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1563_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1563_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext189_1240 : std_logic_vector(31 downto 0);
    signal sext_1296 : std_logic_vector(31 downto 0);
    signal shl_1255 : std_logic_vector(31 downto 0);
    signal shr130_1524 : std_logic_vector(31 downto 0);
    signal shr135_1549 : std_logic_vector(31 downto 0);
    signal shr_1441 : std_logic_vector(31 downto 0);
    signal sub110_1480 : std_logic_vector(31 downto 0);
    signal sub_1470 : std_logic_vector(31 downto 0);
    signal tmp133_1540 : std_logic_vector(63 downto 0);
    signal type_cast_1203_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1238_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1243_wire : std_logic_vector(31 downto 0);
    signal type_cast_1246_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1253_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1268_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1289_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1299_wire : std_logic_vector(31 downto 0);
    signal type_cast_1302_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1312_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1314_wire : std_logic_vector(15 downto 0);
    signal type_cast_1318_wire : std_logic_vector(15 downto 0);
    signal type_cast_1321_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1325_wire : std_logic_vector(15 downto 0);
    signal type_cast_1327_wire : std_logic_vector(15 downto 0);
    signal type_cast_1331_wire : std_logic_vector(31 downto 0);
    signal type_cast_1336_wire : std_logic_vector(31 downto 0);
    signal type_cast_1338_wire : std_logic_vector(31 downto 0);
    signal type_cast_1344_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1349_wire : std_logic_vector(31 downto 0);
    signal type_cast_1351_wire : std_logic_vector(31 downto 0);
    signal type_cast_1368_wire : std_logic_vector(31 downto 0);
    signal type_cast_1373_wire : std_logic_vector(31 downto 0);
    signal type_cast_1375_wire : std_logic_vector(31 downto 0);
    signal type_cast_1381_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1386_wire : std_logic_vector(31 downto 0);
    signal type_cast_1388_wire : std_logic_vector(31 downto 0);
    signal type_cast_1405_wire : std_logic_vector(31 downto 0);
    signal type_cast_1410_wire : std_logic_vector(31 downto 0);
    signal type_cast_1435_wire : std_logic_vector(31 downto 0);
    signal type_cast_1438_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1444_wire : std_logic_vector(63 downto 0);
    signal type_cast_1457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1463_wire : std_logic_vector(31 downto 0);
    signal type_cast_1518_wire : std_logic_vector(31 downto 0);
    signal type_cast_1521_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1527_wire : std_logic_vector(63 downto 0);
    signal type_cast_1543_wire : std_logic_vector(31 downto 0);
    signal type_cast_1546_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1552_wire : std_logic_vector(63 downto 0);
    signal type_cast_1570_wire : std_logic_vector(31 downto 0);
    signal type_cast_1576_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1581_wire : std_logic_vector(31 downto 0);
    signal type_cast_1583_wire : std_logic_vector(31 downto 0);
    signal type_cast_1596_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1604_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1609_wire : std_logic_vector(31 downto 0);
    signal type_cast_1634_wire : std_logic_vector(31 downto 0);
    signal type_cast_1653_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1655_wire : std_logic_vector(15 downto 0);
    signal type_cast_1659_wire : std_logic_vector(15 downto 0);
    signal type_cast_1661_wire : std_logic_vector(15 downto 0);
    signal type_cast_1665_wire : std_logic_vector(15 downto 0);
    signal type_cast_1667_wire : std_logic_vector(15 downto 0);
    signal type_cast_1674_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_1451_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1451_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1451_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1451_resized_base_address <= "00000000000000";
    array_obj_ref_1534_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1534_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1534_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1534_resized_base_address <= "00000000000000";
    array_obj_ref_1559_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1559_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1559_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1559_resized_base_address <= "00000000000000";
    ptr_deref_1455_word_offset_0 <= "00000000000000";
    ptr_deref_1539_word_offset_0 <= "00000000000000";
    ptr_deref_1563_word_offset_0 <= "00000000000000";
    type_cast_1203_wire_constant <= "0000000000000001";
    type_cast_1238_wire_constant <= "00000000000000000000000000010000";
    type_cast_1246_wire_constant <= "00000000000000000000000000010000";
    type_cast_1253_wire_constant <= "00000000000000000000000000000001";
    type_cast_1268_wire_constant <= "00000000000000000000000000000001";
    type_cast_1289_wire_constant <= "00000000000000000000000000010000";
    type_cast_1302_wire_constant <= "00000000000000000000000000010000";
    type_cast_1312_wire_constant <= "0000000000000000";
    type_cast_1321_wire_constant <= "0000000000000000";
    type_cast_1344_wire_constant <= "1";
    type_cast_1381_wire_constant <= "1";
    type_cast_1438_wire_constant <= "00000000000000000000000000000010";
    type_cast_1457_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1521_wire_constant <= "00000000000000000000000000000010";
    type_cast_1546_wire_constant <= "00000000000000000000000000000010";
    type_cast_1576_wire_constant <= "00000000000000000000000000000100";
    type_cast_1596_wire_constant <= "0000000000000100";
    type_cast_1604_wire_constant <= "0000000000000001";
    type_cast_1653_wire_constant <= "0000000000000000";
    type_cast_1674_wire_constant <= "00000001";
    phi_stmt_1308: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1312_wire_constant & type_cast_1314_wire;
      req <= phi_stmt_1308_req_0 & phi_stmt_1308_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1308",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1308_ack_0,
          idata => idata,
          odata => kx_x1_1308,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1308
    phi_stmt_1315: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1318_wire & type_cast_1321_wire_constant;
      req <= phi_stmt_1315_req_0 & phi_stmt_1315_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1315",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1315_ack_0,
          idata => idata,
          odata => ix_x2_1315,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1315
    phi_stmt_1322: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1325_wire & type_cast_1327_wire;
      req <= phi_stmt_1322_req_0 & phi_stmt_1322_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1322",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1322_ack_0,
          idata => idata,
          odata => jx_x1_1322,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1322
    phi_stmt_1649: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1653_wire_constant & type_cast_1655_wire;
      req <= phi_stmt_1649_req_0 & phi_stmt_1649_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1649",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1649_ack_0,
          idata => idata,
          odata => kx_x0x_xph_1649,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1649
    phi_stmt_1656: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1659_wire & type_cast_1661_wire;
      req <= phi_stmt_1656_req_0 & phi_stmt_1656_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1656",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1656_ack_0,
          idata => idata,
          odata => ix_x1x_xph_1656,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1656
    phi_stmt_1662: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1665_wire & type_cast_1667_wire;
      req <= phi_stmt_1662_req_0 & phi_stmt_1662_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1662",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1662_ack_0,
          idata => idata,
          odata => jx_x0x_xph_1662,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1662
    -- flow-through select operator MUX_1630_inst
    jx_x2_1631 <= div_1205 when (cmp160_1616(0) /=  '0') else inc_1606;
    addr_of_1452_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1452_final_reg_req_0;
      addr_of_1452_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1452_final_reg_req_1;
      addr_of_1452_final_reg_ack_1<= rack(0);
      addr_of_1452_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1452_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1451_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1453,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1535_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1535_final_reg_req_0;
      addr_of_1535_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1535_final_reg_req_1;
      addr_of_1535_final_reg_ack_1<= rack(0);
      addr_of_1535_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1535_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1534_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx132_1536,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1560_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1560_final_reg_req_0;
      addr_of_1560_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1560_final_reg_req_1;
      addr_of_1560_final_reg_ack_1<= rack(0);
      addr_of_1560_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1560_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1559_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx137_1561,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1198_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1198_inst_req_0;
      type_cast_1198_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1198_inst_req_1;
      type_cast_1198_inst_ack_1<= rack(0);
      type_cast_1198_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1198_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1199,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1208_inst_req_0;
      type_cast_1208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1208_inst_req_1;
      type_cast_1208_inst_ack_1<= rack(0);
      type_cast_1208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1212_inst_req_0;
      type_cast_1212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1212_inst_req_1;
      type_cast_1212_inst_ack_1<= rack(0);
      type_cast_1212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34_1213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1216_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1216_inst_req_0;
      type_cast_1216_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1216_inst_req_1;
      type_cast_1216_inst_ack_1<= rack(0);
      type_cast_1216_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1216_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_1191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_1217,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1220_inst_req_0;
      type_cast_1220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1220_inst_req_1;
      type_cast_1220_inst_ack_1<= rack(0);
      type_cast_1220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_1188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv40_1221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1229_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1229_inst_req_0;
      type_cast_1229_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1229_inst_req_1;
      type_cast_1229_inst_ack_1<= rack(0);
      type_cast_1229_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1229_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_1230,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1233_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1233_inst_req_0;
      type_cast_1233_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1233_inst_req_1;
      type_cast_1233_inst_ack_1<= rack(0);
      type_cast_1233_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1233_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_1191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_1234,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1243_inst
    process(sext189_1240) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext189_1240(31 downto 0);
      type_cast_1243_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1248_inst
    process(ASHR_i32_i32_1247_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1247_wire(31 downto 0);
      conv87_1249 <= tmp_var; -- 
    end process;
    type_cast_1263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1263_inst_req_0;
      type_cast_1263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1263_inst_req_1;
      type_cast_1263_inst_ack_1<= rack(0);
      type_cast_1263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1264,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1299_inst
    process(sext_1296) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_1296(31 downto 0);
      type_cast_1299_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1304_inst
    process(ASHR_i32_i32_1303_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1303_wire(31 downto 0);
      conv105_1305 <= tmp_var; -- 
    end process;
    type_cast_1314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1314_inst_req_0;
      type_cast_1314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1314_inst_req_1;
      type_cast_1314_inst_ack_1<= rack(0);
      type_cast_1314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_1649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1314_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1318_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1318_inst_req_0;
      type_cast_1318_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1318_inst_req_1;
      type_cast_1318_inst_ack_1<= rack(0);
      type_cast_1318_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1318_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_1656,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1318_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1325_inst_req_0;
      type_cast_1325_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1325_inst_req_1;
      type_cast_1325_inst_ack_1<= rack(0);
      type_cast_1325_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1325_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1205,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1325_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1327_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1327_inst_req_0;
      type_cast_1327_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1327_inst_req_1;
      type_cast_1327_inst_ack_1<= rack(0);
      type_cast_1327_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1327_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_1662,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1327_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1332_inst_req_0;
      type_cast_1332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1332_inst_req_1;
      type_cast_1332_inst_ack_1<= rack(0);
      type_cast_1332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1331_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_1333,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1336_inst
    process(conv47_1333) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv47_1333(31 downto 0);
      type_cast_1336_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1338_inst
    process(conv49_1230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv49_1230(31 downto 0);
      type_cast_1338_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1349_inst
    process(conv47_1333) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv47_1333(31 downto 0);
      type_cast_1349_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1351_inst
    process(add_1280) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_1280(31 downto 0);
      type_cast_1351_wire <= tmp_var; -- 
    end process;
    type_cast_1369_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1369_inst_req_0;
      type_cast_1369_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1369_inst_req_1;
      type_cast_1369_inst_ack_1<= rack(0);
      type_cast_1369_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1369_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1368_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_1370,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1373_inst
    process(conv62_1370) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv62_1370(31 downto 0);
      type_cast_1373_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1375_inst
    process(conv49_1230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv49_1230(31 downto 0);
      type_cast_1375_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1386_inst
    process(conv62_1370) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv62_1370(31 downto 0);
      type_cast_1386_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1388_inst
    process(add74_1285) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add74_1285(31 downto 0);
      type_cast_1388_wire <= tmp_var; -- 
    end process;
    type_cast_1406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1406_inst_req_0;
      type_cast_1406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1406_inst_req_1;
      type_cast_1406_inst_ack_1<= rack(0);
      type_cast_1406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1405_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_1407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1411_inst_req_0;
      type_cast_1411_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1411_inst_req_1;
      type_cast_1411_inst_ack_1<= rack(0);
      type_cast_1411_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1411_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1410_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_1412,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1435_inst
    process(add91_1432) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add91_1432(31 downto 0);
      type_cast_1435_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1440_inst
    process(ASHR_i32_i32_1439_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1439_wire(31 downto 0);
      shr_1441 <= tmp_var; -- 
    end process;
    type_cast_1445_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1445_inst_req_0;
      type_cast_1445_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1445_inst_req_1;
      type_cast_1445_inst_ack_1<= rack(0);
      type_cast_1445_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1445_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1444_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1446,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1464_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1464_inst_req_0;
      type_cast_1464_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1464_inst_req_1;
      type_cast_1464_inst_ack_1<= rack(0);
      type_cast_1464_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1464_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1463_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_1465,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1518_inst
    process(add112_1495) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add112_1495(31 downto 0);
      type_cast_1518_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1523_inst
    process(ASHR_i32_i32_1522_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1522_wire(31 downto 0);
      shr130_1524 <= tmp_var; -- 
    end process;
    type_cast_1528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1528_inst_req_0;
      type_cast_1528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1528_inst_req_1;
      type_cast_1528_inst_ack_1<= rack(0);
      type_cast_1528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1527_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom131_1529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1543_inst
    process(add128_1515) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add128_1515(31 downto 0);
      type_cast_1543_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1548_inst
    process(ASHR_i32_i32_1547_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1547_wire(31 downto 0);
      shr135_1549 <= tmp_var; -- 
    end process;
    type_cast_1553_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1553_inst_req_0;
      type_cast_1553_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1553_inst_req_1;
      type_cast_1553_inst_ack_1<= rack(0);
      type_cast_1553_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1553_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1552_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom136_1554,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1571_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1571_inst_req_0;
      type_cast_1571_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1571_inst_req_1;
      type_cast_1571_inst_ack_1<= rack(0);
      type_cast_1571_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1571_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1570_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv140_1572,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1581_inst
    process(add141_1578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add141_1578(31 downto 0);
      type_cast_1581_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1583_inst
    process(conv32_1209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv32_1209(31 downto 0);
      type_cast_1583_wire <= tmp_var; -- 
    end process;
    type_cast_1610_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1610_inst_req_0;
      type_cast_1610_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1610_inst_req_1;
      type_cast_1610_inst_ack_1<= rack(0);
      type_cast_1610_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1610_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1609_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_1611,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1619_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1619_inst_req_0;
      type_cast_1619_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1619_inst_req_1;
      type_cast_1619_inst_ack_1<= rack(0);
      type_cast_1619_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1619_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp160_1616,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc165_1620,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1635_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1635_inst_req_0;
      type_cast_1635_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1635_inst_req_1;
      type_cast_1635_inst_ack_1<= rack(0);
      type_cast_1635_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1635_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1634_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv168_1636,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1655_inst_req_0;
      type_cast_1655_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1655_inst_req_1;
      type_cast_1655_inst_ack_1<= rack(0);
      type_cast_1655_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add149_1598,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1655_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1659_inst_req_0;
      type_cast_1659_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1659_inst_req_1;
      type_cast_1659_inst_ack_1<= rack(0);
      type_cast_1659_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1659_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc165x_xix_x2_1625,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1659_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1661_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1661_inst_req_0;
      type_cast_1661_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1661_inst_req_1;
      type_cast_1661_inst_ack_1<= rack(0);
      type_cast_1661_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1661_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_1315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1661_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1665_inst_req_0;
      type_cast_1665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1665_inst_req_1;
      type_cast_1665_inst_ack_1<= rack(0);
      type_cast_1665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1665_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_1322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1665_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1667_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1667_inst_req_0;
      type_cast_1667_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1667_inst_req_1;
      type_cast_1667_inst_ack_1<= rack(0);
      type_cast_1667_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1667_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_1631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1667_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1451_index_1_rename
    process(R_idxprom_1450_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1450_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1450_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1451_index_1_resize
    process(idxprom_1446) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1446;
      ov := iv(13 downto 0);
      R_idxprom_1450_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1451_root_address_inst
    process(array_obj_ref_1451_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1451_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1451_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1534_index_1_rename
    process(R_idxprom131_1533_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom131_1533_resized;
      ov(13 downto 0) := iv;
      R_idxprom131_1533_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1534_index_1_resize
    process(idxprom131_1529) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom131_1529;
      ov := iv(13 downto 0);
      R_idxprom131_1533_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1534_root_address_inst
    process(array_obj_ref_1534_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1534_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1534_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1559_index_1_rename
    process(R_idxprom136_1558_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom136_1558_resized;
      ov(13 downto 0) := iv;
      R_idxprom136_1558_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1559_index_1_resize
    process(idxprom136_1554) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom136_1554;
      ov := iv(13 downto 0);
      R_idxprom136_1558_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1559_root_address_inst
    process(array_obj_ref_1559_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1559_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1559_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1455_addr_0
    process(ptr_deref_1455_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1455_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1455_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1455_base_resize
    process(arrayidx_1453) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1453;
      ov := iv(13 downto 0);
      ptr_deref_1455_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1455_gather_scatter
    process(type_cast_1457_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1457_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1455_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1455_root_address_inst
    process(ptr_deref_1455_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1455_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1455_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1539_addr_0
    process(ptr_deref_1539_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1539_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1539_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1539_base_resize
    process(arrayidx132_1536) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx132_1536;
      ov := iv(13 downto 0);
      ptr_deref_1539_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1539_gather_scatter
    process(ptr_deref_1539_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1539_data_0;
      ov(63 downto 0) := iv;
      tmp133_1540 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1539_root_address_inst
    process(ptr_deref_1539_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1539_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1539_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1563_addr_0
    process(ptr_deref_1563_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1563_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1563_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1563_base_resize
    process(arrayidx137_1561) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx137_1561;
      ov := iv(13 downto 0);
      ptr_deref_1563_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1563_gather_scatter
    process(tmp133_1540) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp133_1540;
      ov(63 downto 0) := iv;
      ptr_deref_1563_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1563_root_address_inst
    process(ptr_deref_1563_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1563_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1563_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1359_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_1358;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1359_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1359_branch_req_0,
          ack0 => if_stmt_1359_branch_ack_0,
          ack1 => if_stmt_1359_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1396_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond190_1395;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1396_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1396_branch_req_0,
          ack0 => if_stmt_1396_branch_ack_0,
          ack1 => if_stmt_1396_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1586_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp144_1585;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1586_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1586_branch_req_0,
          ack0 => if_stmt_1586_branch_ack_0,
          ack1 => if_stmt_1586_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1642_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp176_1641;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1642_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1642_branch_req_0,
          ack0 => if_stmt_1642_branch_ack_0,
          ack1 => if_stmt_1642_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1597_inst
    process(kx_x1_1308) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_1308, type_cast_1596_wire_constant, tmp_var);
      add149_1598 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1605_inst
    process(jx_x1_1322) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_1322, type_cast_1604_wire_constant, tmp_var);
      inc_1606 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1624_inst
    process(inc165_1620, ix_x2_1315) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc165_1620, ix_x2_1315, tmp_var);
      inc165x_xix_x2_1625 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1259_inst
    process(shl_1255, conv34_1213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_1255, conv34_1213, tmp_var);
      add159_1260 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1274_inst
    process(shl_1255, div171_1270) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_1255, div171_1270, tmp_var);
      add175_1275 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1279_inst
    process(conv49_1230, div171_1270) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv49_1230, div171_1270, tmp_var);
      add_1280 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1284_inst
    process(conv49_1230, conv34_1213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv49_1230, conv34_1213, tmp_var);
      add74_1285 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1426_inst
    process(mul90_1422, conv79_1407) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul90_1422, conv79_1407, tmp_var);
      add85_1427 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1431_inst
    process(add85_1427, mul84_1417) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add85_1427, mul84_1417, tmp_var);
      add91_1432 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1489_inst
    process(mul111_1485, conv95_1465) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul111_1485, conv95_1465, tmp_var);
      add103_1490 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1494_inst
    process(add103_1490, mul102_1475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add103_1490, mul102_1475, tmp_var);
      add112_1495 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1509_inst
    process(mul127_1505, conv95_1465) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul127_1505, conv95_1465, tmp_var);
      add122_1510 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1514_inst
    process(add122_1510, mul121_1500) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add122_1510, mul121_1500, tmp_var);
      add128_1515 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1577_inst
    process(conv140_1572) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv140_1572, type_cast_1576_wire_constant, tmp_var);
      add141_1578 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1357_inst
    process(cmpx_xnot_1346, cmp58_1353) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_1346, cmp58_1353, tmp_var);
      orx_xcond_1358 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1394_inst
    process(cmp65x_xnot_1383, cmp75_1390) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp65x_xnot_1383, cmp75_1390, tmp_var);
      orx_xcond190_1395 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1247_inst
    process(type_cast_1243_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1243_wire, type_cast_1246_wire_constant, tmp_var);
      ASHR_i32_i32_1247_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1303_inst
    process(type_cast_1299_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1299_wire, type_cast_1302_wire_constant, tmp_var);
      ASHR_i32_i32_1303_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1439_inst
    process(type_cast_1435_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1435_wire, type_cast_1438_wire_constant, tmp_var);
      ASHR_i32_i32_1439_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1522_inst
    process(type_cast_1518_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1518_wire, type_cast_1521_wire_constant, tmp_var);
      ASHR_i32_i32_1522_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1547_inst
    process(type_cast_1543_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1543_wire, type_cast_1546_wire_constant, tmp_var);
      ASHR_i32_i32_1547_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1615_inst
    process(conv154_1611, add159_1260) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv154_1611, add159_1260, tmp_var);
      cmp160_1616 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1640_inst
    process(conv168_1636, add175_1275) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv168_1636, add175_1275, tmp_var);
      cmp176_1641 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1204_inst
    process(conv_1199) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv_1199, type_cast_1203_wire_constant, tmp_var);
      div_1205 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1269_inst
    process(conv170_1264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv170_1264, type_cast_1268_wire_constant, tmp_var);
      div171_1270 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1225_inst
    process(conv38_1217, conv40_1221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv38_1217, conv40_1221, tmp_var);
      mul41_1226 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1295_inst
    process(mul_1291, conv32_1209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1291, conv32_1209, tmp_var);
      sext_1296 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1416_inst
    process(conv83_1412, conv81_1234) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv83_1412, conv81_1234, tmp_var);
      mul84_1417 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1421_inst
    process(conv47_1333, conv87_1249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv47_1333, conv87_1249, tmp_var);
      mul90_1422 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1474_inst
    process(sub_1470, conv32_1209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_1470, conv32_1209, tmp_var);
      mul102_1475 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1484_inst
    process(sub110_1480, conv105_1305) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub110_1480, conv105_1305, tmp_var);
      mul111_1485 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1499_inst
    process(conv62_1370, conv81_1234) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv62_1370, conv81_1234, tmp_var);
      mul121_1500 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1504_inst
    process(conv47_1333, conv87_1249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv47_1333, conv87_1249, tmp_var);
      mul127_1505 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1239_inst
    process(mul41_1226) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul41_1226, type_cast_1238_wire_constant, tmp_var);
      sext189_1240 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1254_inst
    process(conv49_1230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_1230, type_cast_1253_wire_constant, tmp_var);
      shl_1255 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1290_inst
    process(conv34_1213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv34_1213, type_cast_1289_wire_constant, tmp_var);
      mul_1291 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1339_inst
    process(type_cast_1336_wire, type_cast_1338_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1336_wire, type_cast_1338_wire, tmp_var);
      cmp_1340 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1352_inst
    process(type_cast_1349_wire, type_cast_1351_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1349_wire, type_cast_1351_wire, tmp_var);
      cmp58_1353 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1376_inst
    process(type_cast_1373_wire, type_cast_1375_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1373_wire, type_cast_1375_wire, tmp_var);
      cmp65_1377 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1389_inst
    process(type_cast_1386_wire, type_cast_1388_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1386_wire, type_cast_1388_wire, tmp_var);
      cmp75_1390 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1584_inst
    process(type_cast_1581_wire, type_cast_1583_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1581_wire, type_cast_1583_wire, tmp_var);
      cmp144_1585 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1469_inst
    process(conv62_1370, conv49_1230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv62_1370, conv49_1230, tmp_var);
      sub_1470 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1479_inst
    process(conv47_1333, conv49_1230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv47_1333, conv49_1230, tmp_var);
      sub110_1480 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1345_inst
    process(cmp_1340) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_1340, type_cast_1344_wire_constant, tmp_var);
      cmpx_xnot_1346 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1382_inst
    process(cmp65_1377) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp65_1377, type_cast_1381_wire_constant, tmp_var);
      cmp65x_xnot_1383 <= tmp_var; --
    end process;
    -- shared split operator group (45) : array_obj_ref_1451_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1450_scaled;
      array_obj_ref_1451_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1451_index_offset_req_0;
      array_obj_ref_1451_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1451_index_offset_req_1;
      array_obj_ref_1451_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : array_obj_ref_1534_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom131_1533_scaled;
      array_obj_ref_1534_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1534_index_offset_req_0;
      array_obj_ref_1534_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1534_index_offset_req_1;
      array_obj_ref_1534_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_1559_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom136_1558_scaled;
      array_obj_ref_1559_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1559_index_offset_req_0;
      array_obj_ref_1559_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1559_index_offset_req_1;
      array_obj_ref_1559_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- unary operator type_cast_1331_inst
    process(ix_x2_1315) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_1315, tmp_var);
      type_cast_1331_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1368_inst
    process(jx_x1_1322) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1322, tmp_var);
      type_cast_1368_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1405_inst
    process(kx_x1_1308) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1308, tmp_var);
      type_cast_1405_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1410_inst
    process(jx_x1_1322) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1322, tmp_var);
      type_cast_1410_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1444_inst
    process(shr_1441) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1441, tmp_var);
      type_cast_1444_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1463_inst
    process(kx_x1_1308) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1308, tmp_var);
      type_cast_1463_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1527_inst
    process(shr130_1524) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr130_1524, tmp_var);
      type_cast_1527_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1552_inst
    process(shr135_1549) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr135_1549, tmp_var);
      type_cast_1552_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1570_inst
    process(kx_x1_1308) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1308, tmp_var);
      type_cast_1570_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1609_inst
    process(inc_1606) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1606, tmp_var);
      type_cast_1609_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1634_inst
    process(inc165x_xix_x2_1625) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc165x_xix_x2_1625, tmp_var);
      type_cast_1634_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1539_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1539_load_0_req_0;
      ptr_deref_1539_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1539_load_0_req_1;
      ptr_deref_1539_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1539_word_address_0;
      ptr_deref_1539_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1455_store_0 ptr_deref_1563_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1455_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1563_store_0_req_0;
      ptr_deref_1455_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1563_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1455_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1563_store_0_req_1;
      ptr_deref_1455_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1563_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1455_word_address_0 & ptr_deref_1563_word_address_0;
      data_in <= ptr_deref_1455_data_0 & ptr_deref_1563_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_starting_1193_inst RPIPE_Block1_starting_1190_inst RPIPE_Block1_starting_1187_inst RPIPE_Block1_starting_1184_inst RPIPE_Block1_starting_1181_inst RPIPE_Block1_starting_1178_inst RPIPE_Block1_starting_1175_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block1_starting_1193_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_starting_1190_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_starting_1187_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_starting_1184_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_starting_1181_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_starting_1178_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_starting_1175_inst_req_0;
      RPIPE_Block1_starting_1193_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_starting_1190_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_starting_1187_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_starting_1184_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_starting_1181_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_starting_1178_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_starting_1175_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block1_starting_1193_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_starting_1190_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_starting_1187_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_starting_1184_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_starting_1181_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_starting_1178_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_starting_1175_inst_req_1;
      RPIPE_Block1_starting_1193_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_starting_1190_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_starting_1187_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_starting_1184_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_starting_1181_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_starting_1178_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_starting_1175_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call6_1194 <= data_out(55 downto 48);
      call5_1191 <= data_out(47 downto 40);
      call4_1188 <= data_out(39 downto 32);
      call3_1185 <= data_out(31 downto 24);
      call2_1182 <= data_out(23 downto 16);
      call1_1179 <= data_out(15 downto 8);
      call_1176 <= data_out(7 downto 0);
      Block1_starting_read_0_gI: SplitGuardInterface generic map(name => "Block1_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block1_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_starting_pipe_read_req(0),
          oack => Block1_starting_pipe_read_ack(0),
          odata => Block1_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_complete_1672_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_complete_1672_inst_req_0;
      WPIPE_Block1_complete_1672_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_complete_1672_inst_req_1;
      WPIPE_Block1_complete_1672_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1674_wire_constant;
      Block1_complete_write_0_gI: SplitGuardInterface generic map(name => "Block1_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_complete_pipe_write_req(0),
          oack => Block1_complete_pipe_write_ack(0),
          odata => Block1_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_B_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_C is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block2_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_C;
architecture zeropad3D_C_arch of zeropad3D_C is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_C_CP_4296_start: Boolean;
  signal zeropad3D_C_CP_4296_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_Block2_complete_2181_inst_ack_1 : boolean;
  signal array_obj_ref_2067_index_offset_req_0 : boolean;
  signal type_cast_2170_inst_req_0 : boolean;
  signal type_cast_2127_inst_req_0 : boolean;
  signal WPIPE_Block2_complete_2181_inst_req_1 : boolean;
  signal array_obj_ref_2067_index_offset_req_1 : boolean;
  signal type_cast_2127_inst_ack_0 : boolean;
  signal type_cast_1835_inst_ack_0 : boolean;
  signal type_cast_1835_inst_req_0 : boolean;
  signal array_obj_ref_2067_index_offset_ack_0 : boolean;
  signal array_obj_ref_2067_index_offset_ack_1 : boolean;
  signal ptr_deref_2071_store_0_req_1 : boolean;
  signal RPIPE_Block2_starting_1683_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1683_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1683_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1683_inst_ack_1 : boolean;
  signal type_cast_2161_inst_req_0 : boolean;
  signal type_cast_2161_inst_ack_0 : boolean;
  signal phi_stmt_2158_req_1 : boolean;
  signal type_cast_2176_inst_ack_1 : boolean;
  signal type_cast_2127_inst_req_1 : boolean;
  signal phi_stmt_2158_req_0 : boolean;
  signal type_cast_2176_inst_req_1 : boolean;
  signal type_cast_1819_inst_req_0 : boolean;
  signal type_cast_1819_inst_ack_0 : boolean;
  signal type_cast_2118_inst_req_0 : boolean;
  signal type_cast_2161_inst_req_1 : boolean;
  signal type_cast_2161_inst_ack_1 : boolean;
  signal type_cast_2176_inst_ack_0 : boolean;
  signal type_cast_2170_inst_ack_0 : boolean;
  signal phi_stmt_2171_req_1 : boolean;
  signal type_cast_2127_inst_ack_1 : boolean;
  signal phi_stmt_2165_req_1 : boolean;
  signal type_cast_1835_inst_req_1 : boolean;
  signal type_cast_1819_inst_req_1 : boolean;
  signal type_cast_2170_inst_req_1 : boolean;
  signal type_cast_1819_inst_ack_1 : boolean;
  signal phi_stmt_1816_req_0 : boolean;
  signal phi_stmt_1829_req_0 : boolean;
  signal type_cast_2170_inst_ack_1 : boolean;
  signal type_cast_1835_inst_ack_1 : boolean;
  signal phi_stmt_1829_req_1 : boolean;
  signal type_cast_2144_inst_req_0 : boolean;
  signal type_cast_2144_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1686_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1686_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1686_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1686_inst_ack_1 : boolean;
  signal RPIPE_Block2_starting_1689_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1689_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1689_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1689_inst_ack_1 : boolean;
  signal RPIPE_Block2_starting_1692_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1692_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1692_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1692_inst_ack_1 : boolean;
  signal RPIPE_Block2_starting_1695_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1695_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1695_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1695_inst_ack_1 : boolean;
  signal RPIPE_Block2_starting_1698_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1698_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1698_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1698_inst_ack_1 : boolean;
  signal RPIPE_Block2_starting_1701_inst_req_0 : boolean;
  signal RPIPE_Block2_starting_1701_inst_ack_0 : boolean;
  signal RPIPE_Block2_starting_1701_inst_req_1 : boolean;
  signal RPIPE_Block2_starting_1701_inst_ack_1 : boolean;
  signal type_cast_1706_inst_req_0 : boolean;
  signal type_cast_1706_inst_ack_0 : boolean;
  signal type_cast_1706_inst_req_1 : boolean;
  signal type_cast_1706_inst_ack_1 : boolean;
  signal type_cast_1716_inst_req_0 : boolean;
  signal type_cast_1716_inst_ack_0 : boolean;
  signal type_cast_1716_inst_req_1 : boolean;
  signal type_cast_1716_inst_ack_1 : boolean;
  signal type_cast_1720_inst_req_0 : boolean;
  signal type_cast_1720_inst_ack_0 : boolean;
  signal type_cast_1720_inst_req_1 : boolean;
  signal type_cast_1720_inst_ack_1 : boolean;
  signal type_cast_1724_inst_req_0 : boolean;
  signal type_cast_1724_inst_ack_0 : boolean;
  signal type_cast_1724_inst_req_1 : boolean;
  signal type_cast_1724_inst_ack_1 : boolean;
  signal type_cast_1728_inst_req_0 : boolean;
  signal type_cast_1728_inst_ack_0 : boolean;
  signal type_cast_1728_inst_req_1 : boolean;
  signal type_cast_1728_inst_ack_1 : boolean;
  signal type_cast_1737_inst_req_0 : boolean;
  signal type_cast_1737_inst_ack_0 : boolean;
  signal type_cast_1737_inst_req_1 : boolean;
  signal type_cast_1737_inst_ack_1 : boolean;
  signal type_cast_1741_inst_req_0 : boolean;
  signal type_cast_1741_inst_ack_0 : boolean;
  signal type_cast_1741_inst_req_1 : boolean;
  signal type_cast_1741_inst_ack_1 : boolean;
  signal type_cast_1777_inst_req_0 : boolean;
  signal type_cast_1777_inst_ack_0 : boolean;
  signal type_cast_1777_inst_req_1 : boolean;
  signal type_cast_1777_inst_ack_1 : boolean;
  signal type_cast_1840_inst_req_0 : boolean;
  signal type_cast_1840_inst_ack_0 : boolean;
  signal type_cast_1840_inst_req_1 : boolean;
  signal type_cast_1840_inst_ack_1 : boolean;
  signal if_stmt_1867_branch_req_0 : boolean;
  signal if_stmt_1867_branch_ack_1 : boolean;
  signal if_stmt_1867_branch_ack_0 : boolean;
  signal type_cast_1877_inst_req_0 : boolean;
  signal type_cast_1877_inst_ack_0 : boolean;
  signal type_cast_1877_inst_req_1 : boolean;
  signal type_cast_1877_inst_ack_1 : boolean;
  signal if_stmt_1904_branch_req_0 : boolean;
  signal if_stmt_1904_branch_ack_1 : boolean;
  signal if_stmt_1904_branch_ack_0 : boolean;
  signal type_cast_1914_inst_req_0 : boolean;
  signal type_cast_1914_inst_ack_0 : boolean;
  signal type_cast_1914_inst_req_1 : boolean;
  signal type_cast_1914_inst_ack_1 : boolean;
  signal type_cast_1919_inst_req_0 : boolean;
  signal type_cast_1919_inst_ack_0 : boolean;
  signal type_cast_1919_inst_req_1 : boolean;
  signal type_cast_1919_inst_ack_1 : boolean;
  signal type_cast_1953_inst_req_0 : boolean;
  signal type_cast_1953_inst_ack_0 : boolean;
  signal type_cast_1953_inst_req_1 : boolean;
  signal type_cast_1953_inst_ack_1 : boolean;
  signal addr_of_2068_final_reg_ack_1 : boolean;
  signal addr_of_2068_final_reg_req_1 : boolean;
  signal array_obj_ref_1959_index_offset_req_0 : boolean;
  signal WPIPE_Block2_complete_2181_inst_ack_0 : boolean;
  signal array_obj_ref_1959_index_offset_ack_0 : boolean;
  signal array_obj_ref_1959_index_offset_req_1 : boolean;
  signal WPIPE_Block2_complete_2181_inst_req_0 : boolean;
  signal array_obj_ref_1959_index_offset_ack_1 : boolean;
  signal if_stmt_2094_branch_ack_0 : boolean;
  signal phi_stmt_1829_ack_0 : boolean;
  signal addr_of_1960_final_reg_req_0 : boolean;
  signal addr_of_1960_final_reg_ack_0 : boolean;
  signal type_cast_2118_inst_ack_1 : boolean;
  signal addr_of_1960_final_reg_req_1 : boolean;
  signal addr_of_1960_final_reg_ack_1 : boolean;
  signal type_cast_2176_inst_req_0 : boolean;
  signal phi_stmt_1816_req_1 : boolean;
  signal phi_stmt_1823_req_0 : boolean;
  signal type_cast_1826_inst_ack_1 : boolean;
  signal if_stmt_2094_branch_ack_1 : boolean;
  signal type_cast_2118_inst_req_1 : boolean;
  signal phi_stmt_1823_req_1 : boolean;
  signal ptr_deref_2071_store_0_ack_0 : boolean;
  signal ptr_deref_1963_store_0_req_0 : boolean;
  signal ptr_deref_1963_store_0_ack_0 : boolean;
  signal addr_of_2068_final_reg_ack_0 : boolean;
  signal ptr_deref_2071_store_0_req_0 : boolean;
  signal ptr_deref_1963_store_0_req_1 : boolean;
  signal ptr_deref_1963_store_0_ack_1 : boolean;
  signal if_stmt_2094_branch_req_0 : boolean;
  signal phi_stmt_1823_ack_0 : boolean;
  signal phi_stmt_1816_ack_0 : boolean;
  signal type_cast_1826_inst_req_1 : boolean;
  signal type_cast_1828_inst_ack_1 : boolean;
  signal type_cast_1972_inst_req_0 : boolean;
  signal if_stmt_2151_branch_ack_0 : boolean;
  signal type_cast_1972_inst_ack_0 : boolean;
  signal type_cast_1828_inst_req_1 : boolean;
  signal type_cast_1972_inst_req_1 : boolean;
  signal type_cast_1972_inst_ack_1 : boolean;
  signal if_stmt_2151_branch_ack_1 : boolean;
  signal type_cast_2036_inst_req_0 : boolean;
  signal type_cast_2036_inst_ack_0 : boolean;
  signal type_cast_2036_inst_req_1 : boolean;
  signal type_cast_2036_inst_ack_1 : boolean;
  signal addr_of_2068_final_reg_req_0 : boolean;
  signal type_cast_1826_inst_ack_0 : boolean;
  signal type_cast_1826_inst_req_0 : boolean;
  signal type_cast_1828_inst_ack_0 : boolean;
  signal type_cast_2079_inst_ack_1 : boolean;
  signal type_cast_2118_inst_ack_0 : boolean;
  signal type_cast_2079_inst_req_1 : boolean;
  signal array_obj_ref_2042_index_offset_req_0 : boolean;
  signal array_obj_ref_2042_index_offset_ack_0 : boolean;
  signal array_obj_ref_2042_index_offset_req_1 : boolean;
  signal if_stmt_2151_branch_req_0 : boolean;
  signal array_obj_ref_2042_index_offset_ack_1 : boolean;
  signal type_cast_1828_inst_req_0 : boolean;
  signal addr_of_2043_final_reg_req_0 : boolean;
  signal addr_of_2043_final_reg_ack_0 : boolean;
  signal addr_of_2043_final_reg_req_1 : boolean;
  signal addr_of_2043_final_reg_ack_1 : boolean;
  signal type_cast_2079_inst_ack_0 : boolean;
  signal type_cast_2079_inst_req_0 : boolean;
  signal type_cast_2144_inst_ack_1 : boolean;
  signal type_cast_2144_inst_req_1 : boolean;
  signal ptr_deref_2047_load_0_req_0 : boolean;
  signal ptr_deref_2071_store_0_ack_1 : boolean;
  signal ptr_deref_2047_load_0_ack_0 : boolean;
  signal ptr_deref_2047_load_0_req_1 : boolean;
  signal ptr_deref_2047_load_0_ack_1 : boolean;
  signal type_cast_2061_inst_req_0 : boolean;
  signal type_cast_2061_inst_ack_0 : boolean;
  signal type_cast_2061_inst_req_1 : boolean;
  signal type_cast_2061_inst_ack_1 : boolean;
  signal type_cast_2168_inst_req_0 : boolean;
  signal type_cast_2168_inst_ack_0 : boolean;
  signal type_cast_2168_inst_req_1 : boolean;
  signal type_cast_2168_inst_ack_1 : boolean;
  signal phi_stmt_2165_req_0 : boolean;
  signal type_cast_2174_inst_req_0 : boolean;
  signal type_cast_2174_inst_ack_0 : boolean;
  signal type_cast_2174_inst_req_1 : boolean;
  signal type_cast_2174_inst_ack_1 : boolean;
  signal phi_stmt_2171_req_0 : boolean;
  signal phi_stmt_2158_ack_0 : boolean;
  signal phi_stmt_2165_ack_0 : boolean;
  signal phi_stmt_2171_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_C_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_C_CP_4296_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_C_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_C_CP_4296_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_C_CP_4296_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_C_CP_4296_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_C_CP_4296: Block -- control-path 
    signal zeropad3D_C_CP_4296_elements: BooleanArray(134 downto 0);
    -- 
  begin -- 
    zeropad3D_C_CP_4296_elements(0) <= zeropad3D_C_CP_4296_start;
    zeropad3D_C_CP_4296_symbol <= zeropad3D_C_CP_4296_elements(88);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/$entry
      -- CP-element group 0: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1681/$entry
      -- CP-element group 0: 	 branch_block_stmt_1681/branch_block_stmt_1681__entry__
      -- CP-element group 0: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702__entry__
      -- 
    rr_4362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(0), ack => RPIPE_Block2_starting_1683_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	134 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1: 	98 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	101 
    -- CP-element group 1: 	102 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1681/merge_stmt_2157__exit__
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/$entry
      -- CP-element group 1: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/rr
      -- 
    rr_5198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(1), ack => type_cast_1835_inst_req_0); -- 
    rr_5244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(1), ack => type_cast_1819_inst_req_0); -- 
    cr_5203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(1), ack => type_cast_1835_inst_req_1); -- 
    cr_5249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(1), ack => type_cast_1819_inst_req_1); -- 
    cr_5226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(1), ack => type_cast_1828_inst_req_1); -- 
    rr_5221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(1), ack => type_cast_1828_inst_req_0); -- 
    zeropad3D_C_CP_4296_elements(1) <= zeropad3D_C_CP_4296_elements(134);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_Sample/$exit
      -- 
    ra_4363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1683_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(2)); -- 
    cr_4367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(2), ack => RPIPE_Block2_starting_1683_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1683_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_Sample/rr
      -- 
    ca_4368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1683_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(3)); -- 
    rr_4376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(3), ack => RPIPE_Block2_starting_1686_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_Update/cr
      -- 
    ra_4377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1686_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(4)); -- 
    cr_4381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(4), ack => RPIPE_Block2_starting_1686_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1686_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_Sample/rr
      -- 
    ca_4382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1686_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(5)); -- 
    rr_4390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(5), ack => RPIPE_Block2_starting_1689_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_Update/cr
      -- 
    ra_4391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1689_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(6)); -- 
    cr_4395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(6), ack => RPIPE_Block2_starting_1689_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1689_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_Sample/rr
      -- 
    ca_4396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1689_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(7)); -- 
    rr_4404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(7), ack => RPIPE_Block2_starting_1692_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_Update/cr
      -- 
    ra_4405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1692_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(8)); -- 
    cr_4409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(8), ack => RPIPE_Block2_starting_1692_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1692_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_Sample/rr
      -- 
    ca_4410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1692_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(9)); -- 
    rr_4418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(9), ack => RPIPE_Block2_starting_1695_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_Update/cr
      -- 
    ra_4419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1695_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(10)); -- 
    cr_4423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(10), ack => RPIPE_Block2_starting_1695_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1695_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_Sample/rr
      -- 
    ca_4424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1695_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(11)); -- 
    rr_4432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(11), ack => RPIPE_Block2_starting_1698_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_Update/cr
      -- 
    ra_4433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1698_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(12)); -- 
    cr_4437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(12), ack => RPIPE_Block2_starting_1698_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1698_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_Sample/rr
      -- 
    ca_4438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1698_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(13)); -- 
    rr_4446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(13), ack => RPIPE_Block2_starting_1701_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_Update/cr
      -- 
    ra_4447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1701_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(14)); -- 
    cr_4451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(14), ack => RPIPE_Block2_starting_1701_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	30 
    -- CP-element group 15: 	31 
    -- CP-element group 15:  members (55) 
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/$exit
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702__exit__
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813__entry__
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1684_to_assign_stmt_1702/RPIPE_Block2_starting_1701_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_Update/cr
      -- 
    ca_4452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_starting_1701_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(15)); -- 
    rr_4463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1706_inst_req_0); -- 
    cr_4468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1706_inst_req_1); -- 
    rr_4477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1716_inst_req_0); -- 
    cr_4482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1716_inst_req_1); -- 
    rr_4491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1720_inst_req_0); -- 
    cr_4496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1720_inst_req_1); -- 
    rr_4505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1724_inst_req_0); -- 
    cr_4510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1724_inst_req_1); -- 
    rr_4519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1728_inst_req_0); -- 
    cr_4524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1728_inst_req_1); -- 
    rr_4533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1737_inst_req_0); -- 
    cr_4538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1737_inst_req_1); -- 
    rr_4547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1741_inst_req_0); -- 
    cr_4552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1741_inst_req_1); -- 
    rr_4561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1777_inst_req_0); -- 
    cr_4566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(15), ack => type_cast_1777_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_Sample/ra
      -- 
    ra_4464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1706_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1706_Update/ca
      -- 
    ca_4469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1706_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_Sample/ra
      -- 
    ra_4478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1716_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	32 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1716_Update/ca
      -- 
    ca_4483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1716_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_Sample/ra
      -- 
    ra_4492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1720_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	32 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1720_Update/ca
      -- 
    ca_4497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1720_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_Sample/ra
      -- 
    ra_4506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1724_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	32 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1724_Update/ca
      -- 
    ca_4511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1724_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_Sample/ra
      -- 
    ra_4520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1728_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	32 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1728_Update/ca
      -- 
    ca_4525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1728_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_Sample/ra
      -- 
    ra_4534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1737_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	32 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1737_Update/ca
      -- 
    ca_4539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1737_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_Sample/ra
      -- 
    ra_4548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1741_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1741_Update/ca
      -- 
    ca_4553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1741_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_Sample/ra
      -- 
    ra_4562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1777_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/type_cast_1777_Update/ca
      -- 
    ca_4567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1777_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  place  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: 	19 
    -- CP-element group 32: 	21 
    -- CP-element group 32: 	23 
    -- CP-element group 32: 	25 
    -- CP-element group 32: 	27 
    -- CP-element group 32: 	29 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: 	90 
    -- CP-element group 32: 	91 
    -- CP-element group 32: 	93 
    -- CP-element group 32:  members (16) 
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1829/$entry
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/$entry
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813__exit__
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody
      -- CP-element group 32: 	 branch_block_stmt_1681/assign_stmt_1707_to_assign_stmt_1813/$exit
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1816/$entry
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/$entry
      -- 
    cr_5169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(32), ack => type_cast_1826_inst_req_1); -- 
    rr_5164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(32), ack => type_cast_1826_inst_req_0); -- 
    zeropad3D_C_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(17) & zeropad3D_C_CP_4296_elements(19) & zeropad3D_C_CP_4296_elements(21) & zeropad3D_C_CP_4296_elements(23) & zeropad3D_C_CP_4296_elements(25) & zeropad3D_C_CP_4296_elements(27) & zeropad3D_C_CP_4296_elements(29) & zeropad3D_C_CP_4296_elements(31);
      gj_zeropad3D_C_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	109 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_Sample/ra
      -- 
    ra_4579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1840_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(33)); -- 
    -- CP-element group 34:  branch  transition  place  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	109 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (13) 
      -- CP-element group 34: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866__exit__
      -- CP-element group 34: 	 branch_block_stmt_1681/if_stmt_1867__entry__
      -- CP-element group 34: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/$exit
      -- CP-element group 34: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_1681/if_stmt_1867_dead_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1681/if_stmt_1867_eval_test/$entry
      -- CP-element group 34: 	 branch_block_stmt_1681/if_stmt_1867_eval_test/$exit
      -- CP-element group 34: 	 branch_block_stmt_1681/if_stmt_1867_eval_test/branch_req
      -- CP-element group 34: 	 branch_block_stmt_1681/R_orx_xcond_1868_place
      -- CP-element group 34: 	 branch_block_stmt_1681/if_stmt_1867_if_link/$entry
      -- CP-element group 34: 	 branch_block_stmt_1681/if_stmt_1867_else_link/$entry
      -- 
    ca_4584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1840_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(34)); -- 
    branch_req_4592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(34), ack => if_stmt_1867_branch_req_0); -- 
    -- CP-element group 35:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (18) 
      -- CP-element group 35: 	 branch_block_stmt_1681/whilex_xbody_lorx_xlhsx_xfalse58_PhiReq/$entry
      -- CP-element group 35: 	 branch_block_stmt_1681/whilex_xbody_lorx_xlhsx_xfalse58_PhiReq/$exit
      -- CP-element group 35: 	 branch_block_stmt_1681/merge_stmt_1873_PhiAck/$entry
      -- CP-element group 35: 	 branch_block_stmt_1681/merge_stmt_1873_PhiAck/$exit
      -- CP-element group 35: 	 branch_block_stmt_1681/merge_stmt_1873_PhiAck/dummy
      -- CP-element group 35: 	 branch_block_stmt_1681/merge_stmt_1873_PhiReqMerge
      -- CP-element group 35: 	 branch_block_stmt_1681/merge_stmt_1873__exit__
      -- CP-element group 35: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903__entry__
      -- CP-element group 35: 	 branch_block_stmt_1681/if_stmt_1867_if_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_1681/if_stmt_1867_if_link/if_choice_transition
      -- CP-element group 35: 	 branch_block_stmt_1681/whilex_xbody_lorx_xlhsx_xfalse58
      -- CP-element group 35: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/$entry
      -- CP-element group 35: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_Update/cr
      -- 
    if_choice_transition_4597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1867_branch_ack_1, ack => zeropad3D_C_CP_4296_elements(35)); -- 
    rr_4614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(35), ack => type_cast_1877_inst_req_0); -- 
    cr_4619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(35), ack => type_cast_1877_inst_req_1); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	110 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_1681/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_1681/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 36: 	 branch_block_stmt_1681/if_stmt_1867_else_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_1681/if_stmt_1867_else_link/else_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_1681/whilex_xbody_ifx_xthen
      -- 
    else_choice_transition_4601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1867_branch_ack_0, ack => zeropad3D_C_CP_4296_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_Sample/ra
      -- 
    ra_4615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1877_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(37)); -- 
    -- CP-element group 38:  branch  transition  place  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (13) 
      -- CP-element group 38: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903__exit__
      -- CP-element group 38: 	 branch_block_stmt_1681/if_stmt_1904__entry__
      -- CP-element group 38: 	 branch_block_stmt_1681/if_stmt_1904_else_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/$exit
      -- CP-element group 38: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1681/assign_stmt_1878_to_assign_stmt_1903/type_cast_1877_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1681/if_stmt_1904_dead_link/$entry
      -- CP-element group 38: 	 branch_block_stmt_1681/if_stmt_1904_eval_test/$entry
      -- CP-element group 38: 	 branch_block_stmt_1681/if_stmt_1904_eval_test/$exit
      -- CP-element group 38: 	 branch_block_stmt_1681/if_stmt_1904_eval_test/branch_req
      -- CP-element group 38: 	 branch_block_stmt_1681/R_orx_xcond189_1905_place
      -- CP-element group 38: 	 branch_block_stmt_1681/if_stmt_1904_if_link/$entry
      -- 
    ca_4620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1877_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(38)); -- 
    branch_req_4628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(38), ack => if_stmt_1904_branch_req_0); -- 
    -- CP-element group 39:  fork  transition  place  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	55 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	58 
    -- CP-element group 39: 	62 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	66 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	70 
    -- CP-element group 39: 	73 
    -- CP-element group 39:  members (46) 
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_1681/merge_stmt_1968_PhiReqMerge
      -- CP-element group 39: 	 branch_block_stmt_1681/merge_stmt_1968__exit__
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073__entry__
      -- CP-element group 39: 	 branch_block_stmt_1681/if_stmt_1904_if_link/$exit
      -- CP-element group 39: 	 branch_block_stmt_1681/if_stmt_1904_if_link/if_choice_transition
      -- CP-element group 39: 	 branch_block_stmt_1681/lorx_xlhsx_xfalse58_ifx_xelse
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_complete/req
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/merge_stmt_1968_PhiAck/dummy
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1681/merge_stmt_1968_PhiAck/$exit
      -- CP-element group 39: 	 branch_block_stmt_1681/merge_stmt_1968_PhiAck/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1681/lorx_xlhsx_xfalse58_ifx_xelse_PhiReq/$exit
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_final_index_sum_regn_update_start
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_final_index_sum_regn_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_final_index_sum_regn_Update/req
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_complete/req
      -- CP-element group 39: 	 branch_block_stmt_1681/lorx_xlhsx_xfalse58_ifx_xelse_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/word_access_complete/word_0/cr
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_Update/cr
      -- CP-element group 39: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_update_start_
      -- 
    if_choice_transition_4633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1904_branch_ack_1, ack => zeropad3D_C_CP_4296_elements(39)); -- 
    req_4951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(39), ack => array_obj_ref_2067_index_offset_req_1); -- 
    cr_5016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(39), ack => ptr_deref_2071_store_0_req_1); -- 
    req_4966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(39), ack => addr_of_2068_final_reg_req_1); -- 
    rr_4791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(39), ack => type_cast_1972_inst_req_0); -- 
    cr_4796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(39), ack => type_cast_1972_inst_req_1); -- 
    cr_4810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(39), ack => type_cast_2036_inst_req_1); -- 
    req_4841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(39), ack => array_obj_ref_2042_index_offset_req_1); -- 
    req_4856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(39), ack => addr_of_2043_final_reg_req_1); -- 
    cr_4901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(39), ack => ptr_deref_2047_load_0_req_1); -- 
    cr_4920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(39), ack => type_cast_2061_inst_req_1); -- 
    -- CP-element group 40:  transition  place  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	110 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1681/lorx_xlhsx_xfalse58_ifx_xthen_PhiReq/$entry
      -- CP-element group 40: 	 branch_block_stmt_1681/lorx_xlhsx_xfalse58_ifx_xthen_PhiReq/$exit
      -- CP-element group 40: 	 branch_block_stmt_1681/if_stmt_1904_else_link/$exit
      -- CP-element group 40: 	 branch_block_stmt_1681/if_stmt_1904_else_link/else_choice_transition
      -- CP-element group 40: 	 branch_block_stmt_1681/lorx_xlhsx_xfalse58_ifx_xthen
      -- 
    else_choice_transition_4637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1904_branch_ack_0, ack => zeropad3D_C_CP_4296_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	110 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_Sample/ra
      -- 
    ra_4651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1914_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	110 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_Update/ca
      -- 
    ca_4656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1914_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	110 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_Sample/ra
      -- 
    ra_4665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1919_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	110 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_Update/ca
      -- 
    ca_4670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1919_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_Sample/rr
      -- 
    rr_4678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(45), ack => type_cast_1953_inst_req_0); -- 
    zeropad3D_C_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(42) & zeropad3D_C_CP_4296_elements(44);
      gj_zeropad3D_C_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_Sample/ra
      -- 
    ra_4679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	110 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (16) 
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_resized_1
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_scaled_1
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_computed_1
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_resize_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_resize_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_resize_1/index_resize_req
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_resize_1/index_resize_ack
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_scale_1/$entry
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_scale_1/$exit
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_scale_1/scale_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_index_scale_1/scale_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_final_index_sum_regn_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_final_index_sum_regn_Sample/req
      -- 
    ca_4684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(47)); -- 
    req_4709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(47), ack => array_obj_ref_1959_index_offset_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	54 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_final_index_sum_regn_sample_complete
      -- CP-element group 48: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_final_index_sum_regn_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_final_index_sum_regn_Sample/ack
      -- 
    ack_4710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1959_index_offset_ack_0, ack => zeropad3D_C_CP_4296_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	110 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (11) 
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_offset_calculated
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_final_index_sum_regn_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_final_index_sum_regn_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_request/$entry
      -- CP-element group 49: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_request/req
      -- 
    ack_4715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1959_index_offset_ack_1, ack => zeropad3D_C_CP_4296_elements(49)); -- 
    req_4724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(49), ack => addr_of_1960_final_reg_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_request/$exit
      -- CP-element group 50: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_request/ack
      -- 
    ack_4725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1960_final_reg_ack_0, ack => zeropad3D_C_CP_4296_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	110 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (28) 
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_complete/ack
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_base_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_word_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_base_address_resized
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_base_addr_resize/$entry
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_base_addr_resize/$exit
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_base_addr_resize/base_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_base_addr_resize/base_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_word_addrgen/$entry
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_word_addrgen/$exit
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_word_addrgen/root_register_req
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_word_addrgen/root_register_ack
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/ptr_deref_1963_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/ptr_deref_1963_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/ptr_deref_1963_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/ptr_deref_1963_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/word_access_start/word_0/rr
      -- 
    ack_4730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1960_final_reg_ack_1, ack => zeropad3D_C_CP_4296_elements(51)); -- 
    rr_4768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(51), ack => ptr_deref_1963_store_0_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Sample/word_access_start/word_0/ra
      -- 
    ra_4769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_store_0_ack_0, ack => zeropad3D_C_CP_4296_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	110 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Update/word_access_complete/word_0/ca
      -- 
    ca_4780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1963_store_0_ack_1, ack => zeropad3D_C_CP_4296_elements(53)); -- 
    -- CP-element group 54:  join  transition  place  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: 	48 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	111 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1681/ifx_xthen_ifx_xend_PhiReq/$exit
      -- CP-element group 54: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966__exit__
      -- CP-element group 54: 	 branch_block_stmt_1681/ifx_xthen_ifx_xend
      -- CP-element group 54: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/$exit
      -- CP-element group 54: 	 branch_block_stmt_1681/ifx_xthen_ifx_xend_PhiReq/$entry
      -- 
    zeropad3D_C_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(53) & zeropad3D_C_CP_4296_elements(48);
      gj_zeropad3D_C_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	39 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_Sample/ra
      -- 
    ra_4792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1972_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	65 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_1972_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_Sample/rr
      -- 
    ca_4797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1972_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(56)); -- 
    rr_4805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(56), ack => type_cast_2036_inst_req_0); -- 
    rr_4915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(56), ack => type_cast_2061_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_Sample/ra
      -- 
    ra_4806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2036_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	39 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (16) 
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2036_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_final_index_sum_regn_Sample/req
      -- 
    ca_4811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2036_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(58)); -- 
    req_4836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(58), ack => array_obj_ref_2042_index_offset_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	74 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_final_index_sum_regn_Sample/ack
      -- 
    ack_4837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2042_index_offset_ack_0, ack => zeropad3D_C_CP_4296_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2042_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_request/req
      -- 
    ack_4842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2042_index_offset_ack_1, ack => zeropad3D_C_CP_4296_elements(60)); -- 
    req_4851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(60), ack => addr_of_2043_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_request/ack
      -- 
    ack_4852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2043_final_reg_ack_0, ack => zeropad3D_C_CP_4296_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	39 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (24) 
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2043_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Sample/word_access_start/word_0/rr
      -- 
    ack_4857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2043_final_reg_ack_1, ack => zeropad3D_C_CP_4296_elements(62)); -- 
    rr_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(62), ack => ptr_deref_2047_load_0_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Sample/word_access_start/word_0/ra
      -- 
    ra_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2047_load_0_ack_0, ack => zeropad3D_C_CP_4296_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	71 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/ptr_deref_2047_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/ptr_deref_2047_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/ptr_deref_2047_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2047_Update/ptr_deref_2047_Merge/merge_ack
      -- 
    ca_4902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2047_load_0_ack_1, ack => zeropad3D_C_CP_4296_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	56 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_Sample/ra
      -- 
    ra_4916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	39 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_scale_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_final_index_sum_regn_Sample/req
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_final_index_sum_regn_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_scale_1/scale_rename_req
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_scale_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_scale_1/scale_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_resize_1/index_resize_ack
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_resize_1/index_resize_req
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_resize_1/$exit
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_resize_1/$entry
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/type_cast_2061_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_resized_1
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_scaled_1
      -- CP-element group 66: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_index_computed_1
      -- 
    ca_4921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(66)); -- 
    req_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(66), ack => array_obj_ref_2067_index_offset_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	74 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_final_index_sum_regn_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_final_index_sum_regn_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_final_index_sum_regn_sample_complete
      -- 
    ack_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2067_index_offset_ack_0, ack => zeropad3D_C_CP_4296_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (11) 
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_base_plus_offset/$entry
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_final_index_sum_regn_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_final_index_sum_regn_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_base_plus_offset/$exit
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_base_plus_offset/sum_rename_req
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_base_plus_offset/sum_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_request/$entry
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_request/req
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_root_address_calculated
      -- CP-element group 68: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/array_obj_ref_2067_offset_calculated
      -- 
    ack_4952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2067_index_offset_ack_1, ack => zeropad3D_C_CP_4296_elements(68)); -- 
    req_4961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(68), ack => addr_of_2068_final_reg_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_request/ack
      -- CP-element group 69: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_request/$exit
      -- CP-element group 69: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_sample_completed_
      -- 
    ack_4962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2068_final_reg_ack_0, ack => zeropad3D_C_CP_4296_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	39 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (19) 
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_word_addrgen/root_register_req
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_word_addrgen/$entry
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_base_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_word_addrgen/$exit
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_word_addrgen/root_register_ack
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_word_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_base_address_resized
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_base_addr_resize/$entry
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_complete/ack
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_base_addr_resize/base_resize_ack
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_base_addr_resize/base_resize_req
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_base_addr_resize/$exit
      -- CP-element group 70: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/addr_of_2068_update_completed_
      -- 
    ack_4967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2068_final_reg_ack_1, ack => zeropad3D_C_CP_4296_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	64 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/ptr_deref_2071_Split/$entry
      -- CP-element group 71: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/ptr_deref_2071_Split/$exit
      -- CP-element group 71: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/ptr_deref_2071_Split/split_req
      -- CP-element group 71: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/ptr_deref_2071_Split/split_ack
      -- CP-element group 71: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/word_access_start/$entry
      -- CP-element group 71: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/word_access_start/word_0/rr
      -- CP-element group 71: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/word_access_start/word_0/$entry
      -- 
    rr_5005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(71), ack => ptr_deref_2071_store_0_req_0); -- 
    zeropad3D_C_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(64) & zeropad3D_C_CP_4296_elements(70);
      gj_zeropad3D_C_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/word_access_start/$exit
      -- CP-element group 72: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/word_access_start/word_0/ra
      -- CP-element group 72: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Sample/word_access_start/word_0/$exit
      -- 
    ra_5006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2071_store_0_ack_0, ack => zeropad3D_C_CP_4296_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	39 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Update/word_access_complete/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/ptr_deref_2071_Update/word_access_complete/word_0/ca
      -- 
    ca_5017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2071_store_0_ack_1, ack => zeropad3D_C_CP_4296_elements(73)); -- 
    -- CP-element group 74:  join  transition  place  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	59 
    -- CP-element group 74: 	67 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	111 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073__exit__
      -- CP-element group 74: 	 branch_block_stmt_1681/ifx_xelse_ifx_xend
      -- CP-element group 74: 	 branch_block_stmt_1681/ifx_xelse_ifx_xend_PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_1681/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_1681/assign_stmt_1973_to_assign_stmt_2073/$exit
      -- 
    zeropad3D_C_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(59) & zeropad3D_C_CP_4296_elements(67) & zeropad3D_C_CP_4296_elements(73);
      gj_zeropad3D_C_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	111 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_sample_completed_
      -- 
    ra_5029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2079_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(75)); -- 
    -- CP-element group 76:  branch  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	111 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (13) 
      -- CP-element group 76: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093__exit__
      -- CP-element group 76: 	 branch_block_stmt_1681/if_stmt_2094__entry__
      -- CP-element group 76: 	 branch_block_stmt_1681/if_stmt_2094_else_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_1681/if_stmt_2094_if_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_1681/if_stmt_2094_eval_test/branch_req
      -- CP-element group 76: 	 branch_block_stmt_1681/if_stmt_2094_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_1681/R_cmp143_2095_place
      -- CP-element group 76: 	 branch_block_stmt_1681/if_stmt_2094_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_1681/if_stmt_2094_dead_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/$exit
      -- 
    ca_5034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2079_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(76)); -- 
    branch_req_5042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(76), ack => if_stmt_2094_branch_req_0); -- 
    -- CP-element group 77:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	120 
    -- CP-element group 77: 	121 
    -- CP-element group 77: 	123 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	126 
    -- CP-element group 77: 	127 
    -- CP-element group 77:  members (40) 
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xend_ifx_xthen145
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/assign_stmt_2106__entry__
      -- CP-element group 77: 	 branch_block_stmt_1681/assign_stmt_2106__exit__
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xend_ifx_xthen145_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/merge_stmt_2100_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xend_ifx_xthen145_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_1681/merge_stmt_2100_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/merge_stmt_2100_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_1681/merge_stmt_2100_PhiAck/dummy
      -- CP-element group 77: 	 branch_block_stmt_1681/merge_stmt_2100__exit__
      -- CP-element group 77: 	 branch_block_stmt_1681/assign_stmt_2106/$exit
      -- CP-element group 77: 	 branch_block_stmt_1681/assign_stmt_2106/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/if_stmt_2094_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_1681/if_stmt_2094_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/SplitProtocol/Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2094_branch_ack_1, ack => zeropad3D_C_CP_4296_elements(77)); -- 
    rr_5404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(77), ack => type_cast_2161_inst_req_0); -- 
    cr_5409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(77), ack => type_cast_2161_inst_req_1); -- 
    rr_5427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(77), ack => type_cast_2168_inst_req_0); -- 
    cr_5432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(77), ack => type_cast_2168_inst_req_1); -- 
    rr_5450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(77), ack => type_cast_2174_inst_req_0); -- 
    cr_5455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(77), ack => type_cast_2174_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	84 
    -- CP-element group 78:  members (24) 
      -- CP-element group 78: 	 branch_block_stmt_1681/ifx_xend_ifx_xelse150
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1681/merge_stmt_2108__exit__
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150__entry__
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_1681/merge_stmt_2108_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1681/merge_stmt_2108_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_1681/merge_stmt_2108_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1681/merge_stmt_2108_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1681/ifx_xend_ifx_xelse150_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1681/ifx_xend_ifx_xelse150_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/$entry
      -- CP-element group 78: 	 branch_block_stmt_1681/if_stmt_2094_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_1681/if_stmt_2094_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_Update/cr
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_Update/cr
      -- 
    else_choice_transition_5051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2094_branch_ack_0, ack => zeropad3D_C_CP_4296_elements(78)); -- 
    cr_5086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(78), ack => type_cast_2127_inst_req_1); -- 
    rr_5067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(78), ack => type_cast_2118_inst_req_0); -- 
    cr_5072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(78), ack => type_cast_2118_inst_req_1); -- 
    cr_5100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(78), ack => type_cast_2144_inst_req_1); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_Sample/ra
      -- 
    ra_5068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2118_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2118_Update/$exit
      -- 
    ca_5073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2118_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(80)); -- 
    rr_5081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(80), ack => type_cast_2127_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_sample_completed_
      -- 
    ra_5082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2127_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2127_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_Sample/rr
      -- 
    ca_5087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2127_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(82)); -- 
    rr_5095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(82), ack => type_cast_2144_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_Sample/ra
      -- 
    ra_5096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2144_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(83)); -- 
    -- CP-element group 84:  branch  transition  place  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	78 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (13) 
      -- CP-element group 84: 	 branch_block_stmt_1681/R_cmp175_2152_place
      -- CP-element group 84: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150__exit__
      -- CP-element group 84: 	 branch_block_stmt_1681/if_stmt_2151__entry__
      -- CP-element group 84: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/$exit
      -- CP-element group 84: 	 branch_block_stmt_1681/if_stmt_2151_else_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_1681/if_stmt_2151_if_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_1681/if_stmt_2151_eval_test/branch_req
      -- CP-element group 84: 	 branch_block_stmt_1681/if_stmt_2151_eval_test/$exit
      -- CP-element group 84: 	 branch_block_stmt_1681/if_stmt_2151_eval_test/$entry
      -- CP-element group 84: 	 branch_block_stmt_1681/if_stmt_2151_dead_link/$entry
      -- CP-element group 84: 	 branch_block_stmt_1681/assign_stmt_2114_to_assign_stmt_2150/type_cast_2144_Update/ca
      -- 
    ca_5101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2144_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(84)); -- 
    branch_req_5109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(84), ack => if_stmt_2151_branch_req_0); -- 
    -- CP-element group 85:  transition  place  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (15) 
      -- CP-element group 85: 	 branch_block_stmt_1681/ifx_xelse150_whilex_xend
      -- CP-element group 85: 	 branch_block_stmt_1681/merge_stmt_2179__exit__
      -- CP-element group 85: 	 branch_block_stmt_1681/assign_stmt_2184__entry__
      -- CP-element group 85: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1681/assign_stmt_2184/$entry
      -- CP-element group 85: 	 branch_block_stmt_1681/if_stmt_2151_if_link/if_choice_transition
      -- CP-element group 85: 	 branch_block_stmt_1681/if_stmt_2151_if_link/$exit
      -- CP-element group 85: 	 branch_block_stmt_1681/ifx_xelse150_whilex_xend_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_1681/ifx_xelse150_whilex_xend_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1681/merge_stmt_2179_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_1681/merge_stmt_2179_PhiAck/$entry
      -- CP-element group 85: 	 branch_block_stmt_1681/merge_stmt_2179_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_1681/merge_stmt_2179_PhiAck/dummy
      -- 
    if_choice_transition_5114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2151_branch_ack_1, ack => zeropad3D_C_CP_4296_elements(85)); -- 
    req_5131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(85), ack => WPIPE_Block2_complete_2181_inst_req_0); -- 
    -- CP-element group 86:  fork  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	112 
    -- CP-element group 86: 	113 
    -- CP-element group 86: 	114 
    -- CP-element group 86: 	116 
    -- CP-element group 86: 	117 
    -- CP-element group 86:  members (22) 
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2158/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1681/if_stmt_2151_else_link/else_choice_transition
      -- CP-element group 86: 	 branch_block_stmt_1681/if_stmt_2151_else_link/$exit
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/SplitProtocol/Sample/$entry
      -- 
    else_choice_transition_5118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2151_branch_ack_0, ack => zeropad3D_C_CP_4296_elements(86)); -- 
    rr_5355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(86), ack => type_cast_2170_inst_req_0); -- 
    cr_5383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(86), ack => type_cast_2176_inst_req_1); -- 
    cr_5360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(86), ack => type_cast_2170_inst_req_1); -- 
    rr_5378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(86), ack => type_cast_2176_inst_req_0); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_Update/req
      -- CP-element group 87: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_sample_completed_
      -- 
    ack_5132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_complete_2181_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(87)); -- 
    req_5136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(87), ack => WPIPE_Block2_complete_2181_inst_req_1); -- 
    -- CP-element group 88:  transition  place  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1681/return__
      -- CP-element group 88: 	 branch_block_stmt_1681/merge_stmt_2186__exit__
      -- CP-element group 88: 	 branch_block_stmt_1681/assign_stmt_2184__exit__
      -- CP-element group 88: 	 $exit
      -- CP-element group 88: 	 branch_block_stmt_1681/$exit
      -- CP-element group 88: 	 branch_block_stmt_1681/branch_block_stmt_1681__exit__
      -- CP-element group 88: 	 branch_block_stmt_1681/assign_stmt_2184/WPIPE_Block2_complete_2181_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_1681/assign_stmt_2184/$exit
      -- CP-element group 88: 	 branch_block_stmt_1681/return___PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_1681/return___PhiReq/$exit
      -- CP-element group 88: 	 branch_block_stmt_1681/merge_stmt_2186_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_1681/merge_stmt_2186_PhiAck/$entry
      -- CP-element group 88: 	 branch_block_stmt_1681/merge_stmt_2186_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_1681/merge_stmt_2186_PhiAck/dummy
      -- 
    ack_5137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_complete_2181_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(88)); -- 
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	94 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1829/$exit
      -- CP-element group 89: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1833_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_req
      -- 
    phi_stmt_1829_req_5148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1829_req_5148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(89), ack => phi_stmt_1829_req_0); -- 
    -- Element group zeropad3D_C_CP_4296_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => zeropad3D_C_CP_4296_elements(32), ack => zeropad3D_C_CP_4296_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	32 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/$exit
      -- 
    ra_5165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	32 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/$exit
      -- 
    ca_5170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/$exit
      -- CP-element group 92: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_req
      -- CP-element group 92: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/$exit
      -- 
    phi_stmt_1823_req_5171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1823_req_5171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(92), ack => phi_stmt_1823_req_0); -- 
    zeropad3D_C_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(90) & zeropad3D_C_CP_4296_elements(91);
      gj_zeropad3D_C_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  output  delay-element  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	32 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_req
      -- CP-element group 93: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1822_konst_delay_trans
      -- CP-element group 93: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/phi_stmt_1816/$exit
      -- 
    phi_stmt_1816_req_5179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1816_req_5179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(93), ack => phi_stmt_1816_req_1); -- 
    -- Element group zeropad3D_C_CP_4296_elements(93) is a control-delay.
    cp_element_93_delay: control_delay_element  generic map(name => " 93_delay", delay_value => 1)  port map(req => zeropad3D_C_CP_4296_elements(32), ack => zeropad3D_C_CP_4296_elements(93), clk => clk, reset =>reset);
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	89 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	105 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_1681/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(89) & zeropad3D_C_CP_4296_elements(92) & zeropad3D_C_CP_4296_elements(93);
      gj_zeropad3D_C_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/SplitProtocol/Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/SplitProtocol/Sample/$exit
      -- 
    ra_5199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1835_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/SplitProtocol/Update/ca
      -- 
    ca_5204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1835_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	104 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/$exit
      -- CP-element group 97: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/$exit
      -- CP-element group 97: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_sources/type_cast_1835/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1829/phi_stmt_1829_req
      -- 
    phi_stmt_1829_req_5205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1829_req_5205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(97), ack => phi_stmt_1829_req_1); -- 
    zeropad3D_C_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_C_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(95) & zeropad3D_C_CP_4296_elements(96);
      gj_zeropad3D_C_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	1 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/$exit
      -- 
    ra_5222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1828_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/ca
      -- CP-element group 99: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/$exit
      -- 
    ca_5227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1828_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/$exit
      -- CP-element group 100: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_req
      -- CP-element group 100: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/$exit
      -- 
    phi_stmt_1823_req_5228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1823_req_5228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(100), ack => phi_stmt_1823_req_1); -- 
    zeropad3D_C_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(98) & zeropad3D_C_CP_4296_elements(99);
      gj_zeropad3D_C_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	1 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Sample/ra
      -- 
    ra_5245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1819_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Update/ca
      -- 
    ca_5250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1819_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/$exit
      -- CP-element group 103: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/$exit
      -- CP-element group 103: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/phi_stmt_1816_req
      -- CP-element group 103: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/phi_stmt_1816/$exit
      -- 
    phi_stmt_1816_req_5251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1816_req_5251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(103), ack => phi_stmt_1816_req_0); -- 
    zeropad3D_C_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(101) & zeropad3D_C_CP_4296_elements(102);
      gj_zeropad3D_C_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	97 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1681/ifx_xend183_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(97) & zeropad3D_C_CP_4296_elements(100) & zeropad3D_C_CP_4296_elements(103);
      gj_zeropad3D_C_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  merge  fork  transition  place  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	94 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1681/merge_stmt_1815_PhiReqMerge
      -- CP-element group 105: 	 branch_block_stmt_1681/merge_stmt_1815_PhiAck/$entry
      -- 
    zeropad3D_C_CP_4296_elements(105) <= OrReduce(zeropad3D_C_CP_4296_elements(94) & zeropad3D_C_CP_4296_elements(104));
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	109 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1681/merge_stmt_1815_PhiAck/phi_stmt_1816_ack
      -- 
    phi_stmt_1816_ack_5256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1816_ack_0, ack => zeropad3D_C_CP_4296_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_1681/merge_stmt_1815_PhiAck/phi_stmt_1823_ack
      -- 
    phi_stmt_1823_ack_5257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1823_ack_0, ack => zeropad3D_C_CP_4296_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1681/merge_stmt_1815_PhiAck/phi_stmt_1829_ack
      -- 
    phi_stmt_1829_ack_5258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1829_ack_0, ack => zeropad3D_C_CP_4296_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  place  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	106 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	33 
    -- CP-element group 109: 	34 
    -- CP-element group 109:  members (10) 
      -- CP-element group 109: 	 branch_block_stmt_1681/merge_stmt_1815__exit__
      -- CP-element group 109: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866__entry__
      -- CP-element group 109: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/$entry
      -- CP-element group 109: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1681/assign_stmt_1841_to_assign_stmt_1866/type_cast_1840_Update/cr
      -- CP-element group 109: 	 branch_block_stmt_1681/merge_stmt_1815_PhiAck/$exit
      -- 
    rr_4578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(109), ack => type_cast_1840_inst_req_0); -- 
    cr_4583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(109), ack => type_cast_1840_inst_req_1); -- 
    zeropad3D_C_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(106) & zeropad3D_C_CP_4296_elements(107) & zeropad3D_C_CP_4296_elements(108);
      gj_zeropad3D_C_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  merge  fork  transition  place  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	36 
    -- CP-element group 110: 	40 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	53 
    -- CP-element group 110: 	42 
    -- CP-element group 110: 	43 
    -- CP-element group 110: 	44 
    -- CP-element group 110: 	41 
    -- CP-element group 110: 	47 
    -- CP-element group 110: 	49 
    -- CP-element group 110: 	51 
    -- CP-element group 110:  members (33) 
      -- CP-element group 110: 	 branch_block_stmt_1681/merge_stmt_1910_PhiReqMerge
      -- CP-element group 110: 	 branch_block_stmt_1681/merge_stmt_1910_PhiAck/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/merge_stmt_1910_PhiAck/$exit
      -- CP-element group 110: 	 branch_block_stmt_1681/merge_stmt_1910__exit__
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966__entry__
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1914_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1919_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/type_cast_1953_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_final_index_sum_regn_update_start
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_final_index_sum_regn_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/array_obj_ref_1959_final_index_sum_regn_Update/req
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/addr_of_1960_complete/req
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Update/word_access_complete/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Update/word_access_complete/word_0/$entry
      -- CP-element group 110: 	 branch_block_stmt_1681/assign_stmt_1915_to_assign_stmt_1966/ptr_deref_1963_Update/word_access_complete/word_0/cr
      -- CP-element group 110: 	 branch_block_stmt_1681/merge_stmt_1910_PhiAck/dummy
      -- 
    rr_4650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(110), ack => type_cast_1914_inst_req_0); -- 
    cr_4655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(110), ack => type_cast_1914_inst_req_1); -- 
    rr_4664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(110), ack => type_cast_1919_inst_req_0); -- 
    cr_4669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(110), ack => type_cast_1919_inst_req_1); -- 
    cr_4683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(110), ack => type_cast_1953_inst_req_1); -- 
    req_4714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(110), ack => array_obj_ref_1959_index_offset_req_1); -- 
    req_4729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(110), ack => addr_of_1960_final_reg_req_1); -- 
    cr_4779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(110), ack => ptr_deref_1963_store_0_req_1); -- 
    zeropad3D_C_CP_4296_elements(110) <= OrReduce(zeropad3D_C_CP_4296_elements(36) & zeropad3D_C_CP_4296_elements(40));
    -- CP-element group 111:  merge  fork  transition  place  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	54 
    -- CP-element group 111: 	74 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	75 
    -- CP-element group 111: 	76 
    -- CP-element group 111:  members (13) 
      -- CP-element group 111: 	 branch_block_stmt_1681/merge_stmt_2075_PhiAck/$entry
      -- CP-element group 111: 	 branch_block_stmt_1681/merge_stmt_2075_PhiAck/$exit
      -- CP-element group 111: 	 branch_block_stmt_1681/merge_stmt_2075_PhiAck/dummy
      -- CP-element group 111: 	 branch_block_stmt_1681/merge_stmt_2075_PhiReqMerge
      -- CP-element group 111: 	 branch_block_stmt_1681/merge_stmt_2075__exit__
      -- CP-element group 111: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093__entry__
      -- CP-element group 111: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/type_cast_2079_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_1681/assign_stmt_2080_to_assign_stmt_2093/$entry
      -- 
    cr_5033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(111), ack => type_cast_2079_inst_req_1); -- 
    rr_5028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(111), ack => type_cast_2079_inst_req_0); -- 
    zeropad3D_C_CP_4296_elements(111) <= OrReduce(zeropad3D_C_CP_4296_elements(54) & zeropad3D_C_CP_4296_elements(74));
    -- CP-element group 112:  transition  output  delay-element  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	86 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	119 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2164_konst_delay_trans
      -- CP-element group 112: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2158/$exit
      -- CP-element group 112: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_req
      -- CP-element group 112: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/$exit
      -- 
    phi_stmt_2158_req_5339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2158_req_5339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(112), ack => phi_stmt_2158_req_1); -- 
    -- Element group zeropad3D_C_CP_4296_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => zeropad3D_C_CP_4296_elements(86), ack => zeropad3D_C_CP_4296_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	86 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/SplitProtocol/Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/SplitProtocol/Sample/$exit
      -- 
    ra_5356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2170_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	86 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/SplitProtocol/Update/ca
      -- 
    ca_5361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2170_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	119 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/$exit
      -- CP-element group 115: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_req
      -- CP-element group 115: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2170/$exit
      -- CP-element group 115: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/$exit
      -- 
    phi_stmt_2165_req_5362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2165_req_5362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(115), ack => phi_stmt_2165_req_1); -- 
    zeropad3D_C_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(113) & zeropad3D_C_CP_4296_elements(114);
      gj_zeropad3D_C_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	86 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/SplitProtocol/Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/SplitProtocol/Sample/$exit
      -- 
    ra_5379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2176_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	86 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/SplitProtocol/Update/ca
      -- CP-element group 117: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/SplitProtocol/Update/$exit
      -- 
    ca_5384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2176_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2176/$exit
      -- CP-element group 118: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/$exit
      -- CP-element group 118: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_req
      -- CP-element group 118: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/$exit
      -- 
    phi_stmt_2171_req_5385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2171_req_5385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(118), ack => phi_stmt_2171_req_1); -- 
    zeropad3D_C_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(116) & zeropad3D_C_CP_4296_elements(117);
      gj_zeropad3D_C_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	112 
    -- CP-element group 119: 	115 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	130 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1681/ifx_xelse150_ifx_xend183_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(112) & zeropad3D_C_CP_4296_elements(115) & zeropad3D_C_CP_4296_elements(118);
      gj_zeropad3D_C_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	77 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/SplitProtocol/Sample/ra
      -- CP-element group 120: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/SplitProtocol/Sample/$exit
      -- 
    ra_5405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2161_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	77 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/SplitProtocol/Update/ca
      -- CP-element group 121: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/SplitProtocol/Update/$exit
      -- 
    ca_5410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2161_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	129 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/type_cast_2161/$exit
      -- CP-element group 122: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/$exit
      -- CP-element group 122: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_req
      -- CP-element group 122: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2158/phi_stmt_2158_sources/$exit
      -- 
    phi_stmt_2158_req_5411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2158_req_5411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(122), ack => phi_stmt_2158_req_0); -- 
    zeropad3D_C_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(120) & zeropad3D_C_CP_4296_elements(121);
      gj_zeropad3D_C_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	77 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/SplitProtocol/Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/SplitProtocol/Sample/ra
      -- 
    ra_5428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2168_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/SplitProtocol/Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/SplitProtocol/Update/ca
      -- 
    ca_5433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2168_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	129 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/$exit
      -- CP-element group 125: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/$exit
      -- CP-element group 125: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/$exit
      -- CP-element group 125: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_sources/type_cast_2168/SplitProtocol/$exit
      -- CP-element group 125: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2165/phi_stmt_2165_req
      -- 
    phi_stmt_2165_req_5434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2165_req_5434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(125), ack => phi_stmt_2165_req_0); -- 
    zeropad3D_C_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(123) & zeropad3D_C_CP_4296_elements(124);
      gj_zeropad3D_C_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	77 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Sample/ra
      -- 
    ra_5451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2174_inst_ack_0, ack => zeropad3D_C_CP_4296_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	77 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Update/ca
      -- 
    ca_5456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2174_inst_ack_1, ack => zeropad3D_C_CP_4296_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/$exit
      -- CP-element group 128: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/$exit
      -- CP-element group 128: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/$exit
      -- CP-element group 128: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/$exit
      -- CP-element group 128: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/phi_stmt_2171/phi_stmt_2171_req
      -- 
    phi_stmt_2171_req_5457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2171_req_5457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_C_CP_4296_elements(128), ack => phi_stmt_2171_req_0); -- 
    zeropad3D_C_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(126) & zeropad3D_C_CP_4296_elements(127);
      gj_zeropad3D_C_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	122 
    -- CP-element group 129: 	125 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1681/ifx_xthen145_ifx_xend183_PhiReq/$exit
      -- 
    zeropad3D_C_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(122) & zeropad3D_C_CP_4296_elements(125) & zeropad3D_C_CP_4296_elements(128);
      gj_zeropad3D_C_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  fork  transition  place  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	119 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	132 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_1681/merge_stmt_2157_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_1681/merge_stmt_2157_PhiAck/$entry
      -- 
    zeropad3D_C_CP_4296_elements(130) <= OrReduce(zeropad3D_C_CP_4296_elements(119) & zeropad3D_C_CP_4296_elements(129));
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	134 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1681/merge_stmt_2157_PhiAck/phi_stmt_2158_ack
      -- 
    phi_stmt_2158_ack_5462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2158_ack_0, ack => zeropad3D_C_CP_4296_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_1681/merge_stmt_2157_PhiAck/phi_stmt_2165_ack
      -- 
    phi_stmt_2165_ack_5463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2165_ack_0, ack => zeropad3D_C_CP_4296_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_1681/merge_stmt_2157_PhiAck/phi_stmt_2171_ack
      -- 
    phi_stmt_2171_ack_5464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2171_ack_0, ack => zeropad3D_C_CP_4296_elements(133)); -- 
    -- CP-element group 134:  join  transition  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	131 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	1 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_1681/merge_stmt_2157_PhiAck/$exit
      -- 
    zeropad3D_C_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_C_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_C_CP_4296_elements(131) & zeropad3D_C_CP_4296_elements(132) & zeropad3D_C_CP_4296_elements(133);
      gj_zeropad3D_C_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_C_CP_4296_elements(134), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1755_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1811_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1947_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2030_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2055_wire : std_logic_vector(31 downto 0);
    signal R_idxprom130_2041_resized : std_logic_vector(13 downto 0);
    signal R_idxprom130_2041_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom135_2066_resized : std_logic_vector(13 downto 0);
    signal R_idxprom135_2066_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1958_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1958_scaled : std_logic_vector(13 downto 0);
    signal add102_1998 : std_logic_vector(31 downto 0);
    signal add111_2003 : std_logic_vector(31 downto 0);
    signal add121_2018 : std_logic_vector(31 downto 0);
    signal add127_2023 : std_logic_vector(31 downto 0);
    signal add140_2086 : std_logic_vector(31 downto 0);
    signal add148_2106 : std_logic_vector(15 downto 0);
    signal add159_1774 : std_logic_vector(31 downto 0);
    signal add174_1783 : std_logic_vector(31 downto 0);
    signal add73_1793 : std_logic_vector(31 downto 0);
    signal add84_1935 : std_logic_vector(31 downto 0);
    signal add90_1940 : std_logic_vector(31 downto 0);
    signal add_1788 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1959_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1959_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1959_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1959_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1959_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1959_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2042_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2042_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2042_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2042_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2042_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2042_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_root_address : std_logic_vector(13 downto 0);
    signal arrayidx131_2044 : std_logic_vector(31 downto 0);
    signal arrayidx136_2069 : std_logic_vector(31 downto 0);
    signal arrayidx_1961 : std_logic_vector(31 downto 0);
    signal call1_1687 : std_logic_vector(7 downto 0);
    signal call2_1690 : std_logic_vector(7 downto 0);
    signal call3_1693 : std_logic_vector(7 downto 0);
    signal call4_1696 : std_logic_vector(7 downto 0);
    signal call5_1699 : std_logic_vector(7 downto 0);
    signal call6_1702 : std_logic_vector(7 downto 0);
    signal call_1684 : std_logic_vector(7 downto 0);
    signal cmp143_2093 : std_logic_vector(0 downto 0);
    signal cmp160_2124 : std_logic_vector(0 downto 0);
    signal cmp175_2150 : std_logic_vector(0 downto 0);
    signal cmp56_1861 : std_logic_vector(0 downto 0);
    signal cmp63_1885 : std_logic_vector(0 downto 0);
    signal cmp63x_xnot_1891 : std_logic_vector(0 downto 0);
    signal cmp74_1898 : std_logic_vector(0 downto 0);
    signal cmp_1848 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_1854 : std_logic_vector(0 downto 0);
    signal conv104_1813 : std_logic_vector(31 downto 0);
    signal conv139_2080 : std_logic_vector(31 downto 0);
    signal conv153_2119 : std_logic_vector(31 downto 0);
    signal conv168_2145 : std_logic_vector(31 downto 0);
    signal conv170_1778 : std_logic_vector(31 downto 0);
    signal conv31_1717 : std_logic_vector(31 downto 0);
    signal conv33_1721 : std_logic_vector(31 downto 0);
    signal conv37_1725 : std_logic_vector(31 downto 0);
    signal conv39_1729 : std_logic_vector(31 downto 0);
    signal conv46_1841 : std_logic_vector(31 downto 0);
    signal conv48_1738 : std_logic_vector(31 downto 0);
    signal conv60_1878 : std_logic_vector(31 downto 0);
    signal conv78_1915 : std_logic_vector(31 downto 0);
    signal conv80_1742 : std_logic_vector(31 downto 0);
    signal conv82_1920 : std_logic_vector(31 downto 0);
    signal conv86_1757 : std_logic_vector(31 downto 0);
    signal conv94_1973 : std_logic_vector(31 downto 0);
    signal conv_1707 : std_logic_vector(15 downto 0);
    signal div156_1763 : std_logic_vector(31 downto 0);
    signal div_1713 : std_logic_vector(15 downto 0);
    signal idxprom130_2037 : std_logic_vector(63 downto 0);
    signal idxprom135_2062 : std_logic_vector(63 downto 0);
    signal idxprom_1954 : std_logic_vector(63 downto 0);
    signal inc165_2128 : std_logic_vector(15 downto 0);
    signal inc165x_xix_x2_2133 : std_logic_vector(15 downto 0);
    signal inc_2114 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_2165 : std_logic_vector(15 downto 0);
    signal ix_x2_1823 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_2171 : std_logic_vector(15 downto 0);
    signal jx_x1_1829 : std_logic_vector(15 downto 0);
    signal jx_x2_2140 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_2158 : std_logic_vector(15 downto 0);
    signal kx_x1_1816 : std_logic_vector(15 downto 0);
    signal mul101_1983 : std_logic_vector(31 downto 0);
    signal mul110_1993 : std_logic_vector(31 downto 0);
    signal mul120_2008 : std_logic_vector(31 downto 0);
    signal mul126_2013 : std_logic_vector(31 downto 0);
    signal mul40_1734 : std_logic_vector(31 downto 0);
    signal mul83_1925 : std_logic_vector(31 downto 0);
    signal mul89_1930 : std_logic_vector(31 downto 0);
    signal mul_1799 : std_logic_vector(31 downto 0);
    signal orx_xcond189_1903 : std_logic_vector(0 downto 0);
    signal orx_xcond_1866 : std_logic_vector(0 downto 0);
    signal ptr_deref_1963_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1963_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1963_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1963_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1963_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1963_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2047_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2047_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2047_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2047_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2047_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2071_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2071_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2071_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2071_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2071_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2071_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext188_1748 : std_logic_vector(31 downto 0);
    signal sext_1804 : std_logic_vector(31 downto 0);
    signal shl_1769 : std_logic_vector(31 downto 0);
    signal shr129_2032 : std_logic_vector(31 downto 0);
    signal shr134_2057 : std_logic_vector(31 downto 0);
    signal shr_1949 : std_logic_vector(31 downto 0);
    signal sub109_1988 : std_logic_vector(31 downto 0);
    signal sub_1978 : std_logic_vector(31 downto 0);
    signal tmp132_2048 : std_logic_vector(63 downto 0);
    signal type_cast_1711_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1746_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1751_wire : std_logic_vector(31 downto 0);
    signal type_cast_1754_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1761_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1767_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1797_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1807_wire : std_logic_vector(31 downto 0);
    signal type_cast_1810_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1819_wire : std_logic_vector(15 downto 0);
    signal type_cast_1822_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1826_wire : std_logic_vector(15 downto 0);
    signal type_cast_1828_wire : std_logic_vector(15 downto 0);
    signal type_cast_1833_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1835_wire : std_logic_vector(15 downto 0);
    signal type_cast_1839_wire : std_logic_vector(31 downto 0);
    signal type_cast_1844_wire : std_logic_vector(31 downto 0);
    signal type_cast_1846_wire : std_logic_vector(31 downto 0);
    signal type_cast_1852_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1857_wire : std_logic_vector(31 downto 0);
    signal type_cast_1859_wire : std_logic_vector(31 downto 0);
    signal type_cast_1876_wire : std_logic_vector(31 downto 0);
    signal type_cast_1881_wire : std_logic_vector(31 downto 0);
    signal type_cast_1883_wire : std_logic_vector(31 downto 0);
    signal type_cast_1889_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1894_wire : std_logic_vector(31 downto 0);
    signal type_cast_1896_wire : std_logic_vector(31 downto 0);
    signal type_cast_1913_wire : std_logic_vector(31 downto 0);
    signal type_cast_1918_wire : std_logic_vector(31 downto 0);
    signal type_cast_1943_wire : std_logic_vector(31 downto 0);
    signal type_cast_1946_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1952_wire : std_logic_vector(63 downto 0);
    signal type_cast_1965_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1971_wire : std_logic_vector(31 downto 0);
    signal type_cast_2026_wire : std_logic_vector(31 downto 0);
    signal type_cast_2029_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2035_wire : std_logic_vector(63 downto 0);
    signal type_cast_2051_wire : std_logic_vector(31 downto 0);
    signal type_cast_2054_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2060_wire : std_logic_vector(63 downto 0);
    signal type_cast_2078_wire : std_logic_vector(31 downto 0);
    signal type_cast_2084_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2089_wire : std_logic_vector(31 downto 0);
    signal type_cast_2091_wire : std_logic_vector(31 downto 0);
    signal type_cast_2104_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2112_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2117_wire : std_logic_vector(31 downto 0);
    signal type_cast_2137_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2143_wire : std_logic_vector(31 downto 0);
    signal type_cast_2161_wire : std_logic_vector(15 downto 0);
    signal type_cast_2164_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2168_wire : std_logic_vector(15 downto 0);
    signal type_cast_2170_wire : std_logic_vector(15 downto 0);
    signal type_cast_2174_wire : std_logic_vector(15 downto 0);
    signal type_cast_2176_wire : std_logic_vector(15 downto 0);
    signal type_cast_2183_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_1959_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1959_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1959_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1959_resized_base_address <= "00000000000000";
    array_obj_ref_2042_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2042_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2042_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2042_resized_base_address <= "00000000000000";
    array_obj_ref_2067_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2067_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2067_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2067_resized_base_address <= "00000000000000";
    ptr_deref_1963_word_offset_0 <= "00000000000000";
    ptr_deref_2047_word_offset_0 <= "00000000000000";
    ptr_deref_2071_word_offset_0 <= "00000000000000";
    type_cast_1711_wire_constant <= "0000000000000001";
    type_cast_1746_wire_constant <= "00000000000000000000000000010000";
    type_cast_1754_wire_constant <= "00000000000000000000000000010000";
    type_cast_1761_wire_constant <= "00000000000000000000000000000001";
    type_cast_1767_wire_constant <= "00000000000000000000000000000001";
    type_cast_1797_wire_constant <= "00000000000000000000000000010000";
    type_cast_1810_wire_constant <= "00000000000000000000000000010000";
    type_cast_1822_wire_constant <= "0000000000000000";
    type_cast_1833_wire_constant <= "0000000000000000";
    type_cast_1852_wire_constant <= "1";
    type_cast_1889_wire_constant <= "1";
    type_cast_1946_wire_constant <= "00000000000000000000000000000010";
    type_cast_1965_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2029_wire_constant <= "00000000000000000000000000000010";
    type_cast_2054_wire_constant <= "00000000000000000000000000000010";
    type_cast_2084_wire_constant <= "00000000000000000000000000000100";
    type_cast_2104_wire_constant <= "0000000000000100";
    type_cast_2112_wire_constant <= "0000000000000001";
    type_cast_2137_wire_constant <= "0000000000000000";
    type_cast_2164_wire_constant <= "0000000000000000";
    type_cast_2183_wire_constant <= "00000001";
    phi_stmt_1816: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1819_wire & type_cast_1822_wire_constant;
      req <= phi_stmt_1816_req_0 & phi_stmt_1816_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1816",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1816_ack_0,
          idata => idata,
          odata => kx_x1_1816,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1816
    phi_stmt_1823: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1826_wire & type_cast_1828_wire;
      req <= phi_stmt_1823_req_0 & phi_stmt_1823_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1823",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1823_ack_0,
          idata => idata,
          odata => ix_x2_1823,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1823
    phi_stmt_1829: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1833_wire_constant & type_cast_1835_wire;
      req <= phi_stmt_1829_req_0 & phi_stmt_1829_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1829",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1829_ack_0,
          idata => idata,
          odata => jx_x1_1829,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1829
    phi_stmt_2158: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2161_wire & type_cast_2164_wire_constant;
      req <= phi_stmt_2158_req_0 & phi_stmt_2158_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2158",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2158_ack_0,
          idata => idata,
          odata => kx_x0x_xph_2158,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2158
    phi_stmt_2165: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2168_wire & type_cast_2170_wire;
      req <= phi_stmt_2165_req_0 & phi_stmt_2165_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2165",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2165_ack_0,
          idata => idata,
          odata => ix_x1x_xph_2165,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2165
    phi_stmt_2171: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2174_wire & type_cast_2176_wire;
      req <= phi_stmt_2171_req_0 & phi_stmt_2171_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2171",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2171_ack_0,
          idata => idata,
          odata => jx_x0x_xph_2171,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2171
    -- flow-through select operator MUX_2139_inst
    jx_x2_2140 <= type_cast_2137_wire_constant when (cmp160_2124(0) /=  '0') else inc_2114;
    addr_of_1960_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1960_final_reg_req_0;
      addr_of_1960_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1960_final_reg_req_1;
      addr_of_1960_final_reg_ack_1<= rack(0);
      addr_of_1960_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1960_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1959_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1961,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2043_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2043_final_reg_req_0;
      addr_of_2043_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2043_final_reg_req_1;
      addr_of_2043_final_reg_ack_1<= rack(0);
      addr_of_2043_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2043_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2042_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx131_2044,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2068_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2068_final_reg_req_0;
      addr_of_2068_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2068_final_reg_req_1;
      addr_of_2068_final_reg_ack_1<= rack(0);
      addr_of_2068_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2068_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2067_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx136_2069,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1706_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1706_inst_req_0;
      type_cast_1706_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1706_inst_req_1;
      type_cast_1706_inst_ack_1<= rack(0);
      type_cast_1706_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1706_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1707,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1716_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1716_inst_req_0;
      type_cast_1716_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1716_inst_req_1;
      type_cast_1716_inst_ack_1<= rack(0);
      type_cast_1716_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1716_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1690,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_1717,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1720_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1720_inst_req_0;
      type_cast_1720_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1720_inst_req_1;
      type_cast_1720_inst_ack_1<= rack(0);
      type_cast_1720_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1720_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1687,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_1721,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1724_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1724_inst_req_0;
      type_cast_1724_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1724_inst_req_1;
      type_cast_1724_inst_ack_1<= rack(0);
      type_cast_1724_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1724_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_1699,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_1725,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1728_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1728_inst_req_0;
      type_cast_1728_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1728_inst_req_1;
      type_cast_1728_inst_ack_1<= rack(0);
      type_cast_1728_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1728_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_1696,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1729,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1737_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1737_inst_req_0;
      type_cast_1737_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1737_inst_req_1;
      type_cast_1737_inst_ack_1<= rack(0);
      type_cast_1737_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1737_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1702,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_1738,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1741_inst_req_0;
      type_cast_1741_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1741_inst_req_1;
      type_cast_1741_inst_ack_1<= rack(0);
      type_cast_1741_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1741_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_1699,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_1742,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1751_inst
    process(sext188_1748) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext188_1748(31 downto 0);
      type_cast_1751_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1756_inst
    process(ASHR_i32_i32_1755_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1755_wire(31 downto 0);
      conv86_1757 <= tmp_var; -- 
    end process;
    type_cast_1777_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1777_inst_req_0;
      type_cast_1777_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1777_inst_req_1;
      type_cast_1777_inst_ack_1<= rack(0);
      type_cast_1777_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1777_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1778,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1807_inst
    process(sext_1804) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_1804(31 downto 0);
      type_cast_1807_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1812_inst
    process(ASHR_i32_i32_1811_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1811_wire(31 downto 0);
      conv104_1813 <= tmp_var; -- 
    end process;
    type_cast_1819_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1819_inst_req_0;
      type_cast_1819_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1819_inst_req_1;
      type_cast_1819_inst_ack_1<= rack(0);
      type_cast_1819_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1819_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_2158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1819_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1826_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1826_inst_req_0;
      type_cast_1826_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1826_inst_req_1;
      type_cast_1826_inst_ack_1<= rack(0);
      type_cast_1826_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1826_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1713,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1826_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1828_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1828_inst_req_0;
      type_cast_1828_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1828_inst_req_1;
      type_cast_1828_inst_ack_1<= rack(0);
      type_cast_1828_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1828_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_2165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1828_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1835_inst_req_0;
      type_cast_1835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1835_inst_req_1;
      type_cast_1835_inst_ack_1<= rack(0);
      type_cast_1835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_2171,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1835_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1840_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1840_inst_req_0;
      type_cast_1840_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1840_inst_req_1;
      type_cast_1840_inst_ack_1<= rack(0);
      type_cast_1840_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1840_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1839_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv46_1841,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1844_inst
    process(conv46_1841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv46_1841(31 downto 0);
      type_cast_1844_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1846_inst
    process(conv48_1738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv48_1738(31 downto 0);
      type_cast_1846_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1857_inst
    process(conv46_1841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv46_1841(31 downto 0);
      type_cast_1857_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1859_inst
    process(add_1788) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_1788(31 downto 0);
      type_cast_1859_wire <= tmp_var; -- 
    end process;
    type_cast_1877_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1877_inst_req_0;
      type_cast_1877_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1877_inst_req_1;
      type_cast_1877_inst_ack_1<= rack(0);
      type_cast_1877_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1877_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1876_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_1878,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1881_inst
    process(conv60_1878) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv60_1878(31 downto 0);
      type_cast_1881_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1883_inst
    process(conv48_1738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv48_1738(31 downto 0);
      type_cast_1883_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1894_inst
    process(conv60_1878) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv60_1878(31 downto 0);
      type_cast_1894_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1896_inst
    process(add73_1793) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add73_1793(31 downto 0);
      type_cast_1896_wire <= tmp_var; -- 
    end process;
    type_cast_1914_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1914_inst_req_0;
      type_cast_1914_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1914_inst_req_1;
      type_cast_1914_inst_ack_1<= rack(0);
      type_cast_1914_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1914_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1913_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_1915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1919_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1919_inst_req_0;
      type_cast_1919_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1919_inst_req_1;
      type_cast_1919_inst_ack_1<= rack(0);
      type_cast_1919_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1919_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1918_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_1920,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1943_inst
    process(add90_1940) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add90_1940(31 downto 0);
      type_cast_1943_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1948_inst
    process(ASHR_i32_i32_1947_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1947_wire(31 downto 0);
      shr_1949 <= tmp_var; -- 
    end process;
    type_cast_1953_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1953_inst_req_0;
      type_cast_1953_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1953_inst_req_1;
      type_cast_1953_inst_ack_1<= rack(0);
      type_cast_1953_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1953_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1952_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1954,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1972_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1972_inst_req_0;
      type_cast_1972_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1972_inst_req_1;
      type_cast_1972_inst_ack_1<= rack(0);
      type_cast_1972_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1972_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1971_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1973,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2026_inst
    process(add111_2003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add111_2003(31 downto 0);
      type_cast_2026_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2031_inst
    process(ASHR_i32_i32_2030_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2030_wire(31 downto 0);
      shr129_2032 <= tmp_var; -- 
    end process;
    type_cast_2036_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2036_inst_req_0;
      type_cast_2036_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2036_inst_req_1;
      type_cast_2036_inst_ack_1<= rack(0);
      type_cast_2036_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2036_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2035_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom130_2037,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2051_inst
    process(add127_2023) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add127_2023(31 downto 0);
      type_cast_2051_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2056_inst
    process(ASHR_i32_i32_2055_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2055_wire(31 downto 0);
      shr134_2057 <= tmp_var; -- 
    end process;
    type_cast_2061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2061_inst_req_0;
      type_cast_2061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2061_inst_req_1;
      type_cast_2061_inst_ack_1<= rack(0);
      type_cast_2061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2060_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom135_2062,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2079_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2079_inst_req_0;
      type_cast_2079_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2079_inst_req_1;
      type_cast_2079_inst_ack_1<= rack(0);
      type_cast_2079_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2079_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2078_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv139_2080,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2089_inst
    process(add140_2086) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add140_2086(31 downto 0);
      type_cast_2089_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2091_inst
    process(conv31_1717) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv31_1717(31 downto 0);
      type_cast_2091_wire <= tmp_var; -- 
    end process;
    type_cast_2118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2118_inst_req_0;
      type_cast_2118_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2118_inst_req_1;
      type_cast_2118_inst_ack_1<= rack(0);
      type_cast_2118_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2118_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2117_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_2119,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2127_inst_req_0;
      type_cast_2127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2127_inst_req_1;
      type_cast_2127_inst_ack_1<= rack(0);
      type_cast_2127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp160_2124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc165_2128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2144_inst_req_0;
      type_cast_2144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2144_inst_req_1;
      type_cast_2144_inst_ack_1<= rack(0);
      type_cast_2144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2143_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv168_2145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2161_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2161_inst_req_0;
      type_cast_2161_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2161_inst_req_1;
      type_cast_2161_inst_ack_1<= rack(0);
      type_cast_2161_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2161_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add148_2106,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2161_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2168_inst_req_0;
      type_cast_2168_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2168_inst_req_1;
      type_cast_2168_inst_ack_1<= rack(0);
      type_cast_2168_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2168_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_1823,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2168_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2170_inst_req_0;
      type_cast_2170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2170_inst_req_1;
      type_cast_2170_inst_ack_1<= rack(0);
      type_cast_2170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc165x_xix_x2_2133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2170_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2174_inst_req_0;
      type_cast_2174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2174_inst_req_1;
      type_cast_2174_inst_ack_1<= rack(0);
      type_cast_2174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_1829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2174_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2176_inst_req_0;
      type_cast_2176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2176_inst_req_1;
      type_cast_2176_inst_ack_1<= rack(0);
      type_cast_2176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_2140,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2176_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1959_index_1_rename
    process(R_idxprom_1958_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1958_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1958_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1959_index_1_resize
    process(idxprom_1954) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1954;
      ov := iv(13 downto 0);
      R_idxprom_1958_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1959_root_address_inst
    process(array_obj_ref_1959_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1959_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1959_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2042_index_1_rename
    process(R_idxprom130_2041_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom130_2041_resized;
      ov(13 downto 0) := iv;
      R_idxprom130_2041_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2042_index_1_resize
    process(idxprom130_2037) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom130_2037;
      ov := iv(13 downto 0);
      R_idxprom130_2041_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2042_root_address_inst
    process(array_obj_ref_2042_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2042_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2042_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2067_index_1_rename
    process(R_idxprom135_2066_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom135_2066_resized;
      ov(13 downto 0) := iv;
      R_idxprom135_2066_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2067_index_1_resize
    process(idxprom135_2062) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom135_2062;
      ov := iv(13 downto 0);
      R_idxprom135_2066_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2067_root_address_inst
    process(array_obj_ref_2067_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2067_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2067_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1963_addr_0
    process(ptr_deref_1963_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1963_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1963_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1963_base_resize
    process(arrayidx_1961) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1961;
      ov := iv(13 downto 0);
      ptr_deref_1963_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1963_gather_scatter
    process(type_cast_1965_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1965_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1963_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1963_root_address_inst
    process(ptr_deref_1963_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1963_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1963_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2047_addr_0
    process(ptr_deref_2047_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2047_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2047_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2047_base_resize
    process(arrayidx131_2044) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx131_2044;
      ov := iv(13 downto 0);
      ptr_deref_2047_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2047_gather_scatter
    process(ptr_deref_2047_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2047_data_0;
      ov(63 downto 0) := iv;
      tmp132_2048 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2047_root_address_inst
    process(ptr_deref_2047_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2047_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2047_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2071_addr_0
    process(ptr_deref_2071_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2071_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2071_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2071_base_resize
    process(arrayidx136_2069) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx136_2069;
      ov := iv(13 downto 0);
      ptr_deref_2071_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2071_gather_scatter
    process(tmp132_2048) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp132_2048;
      ov(63 downto 0) := iv;
      ptr_deref_2071_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2071_root_address_inst
    process(ptr_deref_2071_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2071_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2071_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1867_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_1866;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1867_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1867_branch_req_0,
          ack0 => if_stmt_1867_branch_ack_0,
          ack1 => if_stmt_1867_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1904_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond189_1903;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1904_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1904_branch_req_0,
          ack0 => if_stmt_1904_branch_ack_0,
          ack1 => if_stmt_1904_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2094_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp143_2093;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2094_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2094_branch_req_0,
          ack0 => if_stmt_2094_branch_ack_0,
          ack1 => if_stmt_2094_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2151_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp175_2150;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2151_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2151_branch_req_0,
          ack0 => if_stmt_2151_branch_ack_0,
          ack1 => if_stmt_2151_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2105_inst
    process(kx_x1_1816) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_1816, type_cast_2104_wire_constant, tmp_var);
      add148_2106 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2113_inst
    process(jx_x1_1829) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_1829, type_cast_2112_wire_constant, tmp_var);
      inc_2114 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2132_inst
    process(inc165_2128, ix_x2_1823) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc165_2128, ix_x2_1823, tmp_var);
      inc165x_xix_x2_2133 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1773_inst
    process(shl_1769, div156_1763) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_1769, div156_1763, tmp_var);
      add159_1774 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1782_inst
    process(shl_1769, conv170_1778) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_1769, conv170_1778, tmp_var);
      add174_1783 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1787_inst
    process(conv48_1738, conv170_1778) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv48_1738, conv170_1778, tmp_var);
      add_1788 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1792_inst
    process(conv48_1738, div156_1763) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv48_1738, div156_1763, tmp_var);
      add73_1793 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1934_inst
    process(mul89_1930, conv78_1915) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul89_1930, conv78_1915, tmp_var);
      add84_1935 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1939_inst
    process(add84_1935, mul83_1925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add84_1935, mul83_1925, tmp_var);
      add90_1940 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1997_inst
    process(mul110_1993, conv94_1973) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul110_1993, conv94_1973, tmp_var);
      add102_1998 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2002_inst
    process(add102_1998, mul101_1983) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add102_1998, mul101_1983, tmp_var);
      add111_2003 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2017_inst
    process(mul126_2013, conv94_1973) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul126_2013, conv94_1973, tmp_var);
      add121_2018 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2022_inst
    process(add121_2018, mul120_2008) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add121_2018, mul120_2008, tmp_var);
      add127_2023 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2085_inst
    process(conv139_2080) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv139_2080, type_cast_2084_wire_constant, tmp_var);
      add140_2086 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1865_inst
    process(cmpx_xnot_1854, cmp56_1861) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_1854, cmp56_1861, tmp_var);
      orx_xcond_1866 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1902_inst
    process(cmp63x_xnot_1891, cmp74_1898) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp63x_xnot_1891, cmp74_1898, tmp_var);
      orx_xcond189_1903 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1755_inst
    process(type_cast_1751_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1751_wire, type_cast_1754_wire_constant, tmp_var);
      ASHR_i32_i32_1755_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1811_inst
    process(type_cast_1807_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1807_wire, type_cast_1810_wire_constant, tmp_var);
      ASHR_i32_i32_1811_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1947_inst
    process(type_cast_1943_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1943_wire, type_cast_1946_wire_constant, tmp_var);
      ASHR_i32_i32_1947_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2030_inst
    process(type_cast_2026_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2026_wire, type_cast_2029_wire_constant, tmp_var);
      ASHR_i32_i32_2030_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2055_inst
    process(type_cast_2051_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2051_wire, type_cast_2054_wire_constant, tmp_var);
      ASHR_i32_i32_2055_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2123_inst
    process(conv153_2119, add159_1774) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv153_2119, add159_1774, tmp_var);
      cmp160_2124 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2149_inst
    process(conv168_2145, add174_1783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv168_2145, add174_1783, tmp_var);
      cmp175_2150 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1712_inst
    process(conv_1707) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv_1707, type_cast_1711_wire_constant, tmp_var);
      div_1713 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1762_inst
    process(conv33_1721) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv33_1721, type_cast_1761_wire_constant, tmp_var);
      div156_1763 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1733_inst
    process(conv37_1725, conv39_1729) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv37_1725, conv39_1729, tmp_var);
      mul40_1734 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1803_inst
    process(mul_1799, conv31_1717) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1799, conv31_1717, tmp_var);
      sext_1804 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1924_inst
    process(conv82_1920, conv80_1742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv82_1920, conv80_1742, tmp_var);
      mul83_1925 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1929_inst
    process(conv46_1841, conv86_1757) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_1841, conv86_1757, tmp_var);
      mul89_1930 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1982_inst
    process(sub_1978, conv31_1717) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_1978, conv31_1717, tmp_var);
      mul101_1983 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1992_inst
    process(sub109_1988, conv104_1813) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub109_1988, conv104_1813, tmp_var);
      mul110_1993 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2007_inst
    process(conv60_1878, conv80_1742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv60_1878, conv80_1742, tmp_var);
      mul120_2008 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2012_inst
    process(conv46_1841, conv86_1757) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_1841, conv86_1757, tmp_var);
      mul126_2013 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1747_inst
    process(mul40_1734) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul40_1734, type_cast_1746_wire_constant, tmp_var);
      sext188_1748 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1768_inst
    process(conv48_1738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv48_1738, type_cast_1767_wire_constant, tmp_var);
      shl_1769 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1798_inst
    process(conv33_1721) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv33_1721, type_cast_1797_wire_constant, tmp_var);
      mul_1799 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1847_inst
    process(type_cast_1844_wire, type_cast_1846_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1844_wire, type_cast_1846_wire, tmp_var);
      cmp_1848 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1860_inst
    process(type_cast_1857_wire, type_cast_1859_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1857_wire, type_cast_1859_wire, tmp_var);
      cmp56_1861 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1884_inst
    process(type_cast_1881_wire, type_cast_1883_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1881_wire, type_cast_1883_wire, tmp_var);
      cmp63_1885 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1897_inst
    process(type_cast_1894_wire, type_cast_1896_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1894_wire, type_cast_1896_wire, tmp_var);
      cmp74_1898 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2092_inst
    process(type_cast_2089_wire, type_cast_2091_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2089_wire, type_cast_2091_wire, tmp_var);
      cmp143_2093 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1977_inst
    process(conv60_1878, conv48_1738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv60_1878, conv48_1738, tmp_var);
      sub_1978 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1987_inst
    process(conv46_1841, conv48_1738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv46_1841, conv48_1738, tmp_var);
      sub109_1988 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1853_inst
    process(cmp_1848) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_1848, type_cast_1852_wire_constant, tmp_var);
      cmpx_xnot_1854 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1890_inst
    process(cmp63_1885) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp63_1885, type_cast_1889_wire_constant, tmp_var);
      cmp63x_xnot_1891 <= tmp_var; --
    end process;
    -- shared split operator group (45) : array_obj_ref_1959_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1958_scaled;
      array_obj_ref_1959_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1959_index_offset_req_0;
      array_obj_ref_1959_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1959_index_offset_req_1;
      array_obj_ref_1959_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : array_obj_ref_2042_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom130_2041_scaled;
      array_obj_ref_2042_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2042_index_offset_req_0;
      array_obj_ref_2042_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2042_index_offset_req_1;
      array_obj_ref_2042_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_2067_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom135_2066_scaled;
      array_obj_ref_2067_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2067_index_offset_req_0;
      array_obj_ref_2067_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2067_index_offset_req_1;
      array_obj_ref_2067_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- unary operator type_cast_1839_inst
    process(ix_x2_1823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_1823, tmp_var);
      type_cast_1839_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1876_inst
    process(jx_x1_1829) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1829, tmp_var);
      type_cast_1876_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1913_inst
    process(kx_x1_1816) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1816, tmp_var);
      type_cast_1913_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1918_inst
    process(jx_x1_1829) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_1829, tmp_var);
      type_cast_1918_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1952_inst
    process(shr_1949) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1949, tmp_var);
      type_cast_1952_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1971_inst
    process(kx_x1_1816) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1816, tmp_var);
      type_cast_1971_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2035_inst
    process(shr129_2032) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr129_2032, tmp_var);
      type_cast_2035_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2060_inst
    process(shr134_2057) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr134_2057, tmp_var);
      type_cast_2060_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2078_inst
    process(kx_x1_1816) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_1816, tmp_var);
      type_cast_2078_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2117_inst
    process(inc_2114) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2114, tmp_var);
      type_cast_2117_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2143_inst
    process(inc165x_xix_x2_2133) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc165x_xix_x2_2133, tmp_var);
      type_cast_2143_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2047_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2047_load_0_req_0;
      ptr_deref_2047_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2047_load_0_req_1;
      ptr_deref_2047_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2047_word_address_0;
      ptr_deref_2047_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1963_store_0 ptr_deref_2071_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1963_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2071_store_0_req_0;
      ptr_deref_1963_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2071_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1963_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2071_store_0_req_1;
      ptr_deref_1963_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2071_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1963_word_address_0 & ptr_deref_2071_word_address_0;
      data_in <= ptr_deref_1963_data_0 & ptr_deref_2071_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_starting_1683_inst RPIPE_Block2_starting_1686_inst RPIPE_Block2_starting_1689_inst RPIPE_Block2_starting_1692_inst RPIPE_Block2_starting_1695_inst RPIPE_Block2_starting_1698_inst RPIPE_Block2_starting_1701_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block2_starting_1683_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_starting_1686_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_starting_1689_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_starting_1692_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_starting_1695_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_starting_1698_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_starting_1701_inst_req_0;
      RPIPE_Block2_starting_1683_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_starting_1686_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_starting_1689_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_starting_1692_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_starting_1695_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_starting_1698_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_starting_1701_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block2_starting_1683_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_starting_1686_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_starting_1689_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_starting_1692_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_starting_1695_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_starting_1698_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_starting_1701_inst_req_1;
      RPIPE_Block2_starting_1683_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_starting_1686_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_starting_1689_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_starting_1692_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_starting_1695_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_starting_1698_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_starting_1701_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call_1684 <= data_out(55 downto 48);
      call1_1687 <= data_out(47 downto 40);
      call2_1690 <= data_out(39 downto 32);
      call3_1693 <= data_out(31 downto 24);
      call4_1696 <= data_out(23 downto 16);
      call5_1699 <= data_out(15 downto 8);
      call6_1702 <= data_out(7 downto 0);
      Block2_starting_read_0_gI: SplitGuardInterface generic map(name => "Block2_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block2_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_starting_pipe_read_req(0),
          oack => Block2_starting_pipe_read_ack(0),
          odata => Block2_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_complete_2181_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_complete_2181_inst_req_0;
      WPIPE_Block2_complete_2181_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_complete_2181_inst_req_1;
      WPIPE_Block2_complete_2181_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2183_wire_constant;
      Block2_complete_write_0_gI: SplitGuardInterface generic map(name => "Block2_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_complete_pipe_write_req(0),
          oack => Block2_complete_pipe_write_ack(0),
          odata => Block2_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_C_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block3_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block3_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_D;
architecture zeropad3D_D_arch of zeropad3D_D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_D_CP_5481_start: Boolean;
  signal zeropad3D_D_CP_5481_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_2554_index_offset_req_1 : boolean;
  signal array_obj_ref_2554_index_offset_ack_1 : boolean;
  signal array_obj_ref_2554_index_offset_ack_0 : boolean;
  signal addr_of_2555_final_reg_req_1 : boolean;
  signal ptr_deref_2475_store_0_req_1 : boolean;
  signal addr_of_2555_final_reg_ack_1 : boolean;
  signal ptr_deref_2475_store_0_ack_1 : boolean;
  signal type_cast_2243_inst_req_0 : boolean;
  signal type_cast_2243_inst_ack_0 : boolean;
  signal type_cast_2431_inst_ack_1 : boolean;
  signal type_cast_2260_inst_req_1 : boolean;
  signal type_cast_2352_inst_ack_0 : boolean;
  signal type_cast_2431_inst_req_1 : boolean;
  signal ptr_deref_2475_store_0_ack_0 : boolean;
  signal addr_of_2472_final_reg_req_1 : boolean;
  signal type_cast_2484_inst_req_0 : boolean;
  signal type_cast_2484_inst_ack_0 : boolean;
  signal type_cast_2548_inst_req_1 : boolean;
  signal type_cast_2389_inst_req_1 : boolean;
  signal array_obj_ref_2471_index_offset_req_1 : boolean;
  signal array_obj_ref_2471_index_offset_ack_1 : boolean;
  signal type_cast_2484_inst_req_1 : boolean;
  signal type_cast_2484_inst_ack_1 : boolean;
  signal addr_of_2555_final_reg_req_0 : boolean;
  signal type_cast_2389_inst_ack_1 : boolean;
  signal type_cast_2247_inst_ack_0 : boolean;
  signal ptr_deref_2559_load_0_req_1 : boolean;
  signal array_obj_ref_2554_index_offset_req_0 : boolean;
  signal ptr_deref_2559_load_0_ack_1 : boolean;
  signal ptr_deref_2559_load_0_req_0 : boolean;
  signal type_cast_2548_inst_ack_1 : boolean;
  signal type_cast_2548_inst_req_0 : boolean;
  signal type_cast_2243_inst_req_1 : boolean;
  signal type_cast_2243_inst_ack_1 : boolean;
  signal type_cast_2256_inst_req_1 : boolean;
  signal type_cast_2247_inst_req_1 : boolean;
  signal if_stmt_2416_branch_req_0 : boolean;
  signal type_cast_2352_inst_req_1 : boolean;
  signal type_cast_2352_inst_ack_1 : boolean;
  signal type_cast_2247_inst_ack_1 : boolean;
  signal addr_of_2555_final_reg_ack_0 : boolean;
  signal type_cast_2256_inst_ack_1 : boolean;
  signal type_cast_2260_inst_ack_1 : boolean;
  signal type_cast_2352_inst_req_0 : boolean;
  signal type_cast_2548_inst_ack_0 : boolean;
  signal addr_of_2472_final_reg_ack_1 : boolean;
  signal type_cast_2573_inst_req_0 : boolean;
  signal type_cast_2573_inst_ack_0 : boolean;
  signal type_cast_2573_inst_req_1 : boolean;
  signal type_cast_2573_inst_ack_1 : boolean;
  signal type_cast_2465_inst_ack_1 : boolean;
  signal array_obj_ref_2471_index_offset_ack_0 : boolean;
  signal type_cast_2256_inst_ack_0 : boolean;
  signal type_cast_2260_inst_ack_0 : boolean;
  signal type_cast_2247_inst_req_0 : boolean;
  signal type_cast_2260_inst_req_0 : boolean;
  signal type_cast_2256_inst_req_0 : boolean;
  signal type_cast_2239_inst_ack_1 : boolean;
  signal type_cast_2389_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2192_inst_req_0 : boolean;
  signal type_cast_2389_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2192_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2192_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2192_inst_ack_1 : boolean;
  signal type_cast_2431_inst_ack_0 : boolean;
  signal array_obj_ref_2471_index_offset_req_0 : boolean;
  signal type_cast_2290_inst_ack_1 : boolean;
  signal RPIPE_Block3_starting_2195_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2195_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2195_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2195_inst_ack_1 : boolean;
  signal type_cast_2431_inst_req_0 : boolean;
  signal type_cast_2290_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2198_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2198_inst_ack_0 : boolean;
  signal type_cast_2465_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2198_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2198_inst_ack_1 : boolean;
  signal type_cast_2290_inst_ack_0 : boolean;
  signal type_cast_2290_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2201_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2201_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2201_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2201_inst_ack_1 : boolean;
  signal ptr_deref_2475_store_0_req_0 : boolean;
  signal type_cast_2426_inst_ack_1 : boolean;
  signal type_cast_2426_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2204_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2204_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2204_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2204_inst_ack_1 : boolean;
  signal RPIPE_Block3_starting_2207_inst_req_0 : boolean;
  signal if_stmt_2379_branch_ack_0 : boolean;
  signal RPIPE_Block3_starting_2207_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2207_inst_req_1 : boolean;
  signal RPIPE_Block3_starting_2207_inst_ack_1 : boolean;
  signal type_cast_2426_inst_ack_0 : boolean;
  signal type_cast_2426_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2210_inst_req_0 : boolean;
  signal RPIPE_Block3_starting_2210_inst_ack_0 : boolean;
  signal RPIPE_Block3_starting_2210_inst_req_1 : boolean;
  signal if_stmt_2379_branch_ack_1 : boolean;
  signal RPIPE_Block3_starting_2210_inst_ack_1 : boolean;
  signal type_cast_2215_inst_req_0 : boolean;
  signal type_cast_2215_inst_ack_0 : boolean;
  signal type_cast_2465_inst_ack_0 : boolean;
  signal type_cast_2465_inst_req_0 : boolean;
  signal type_cast_2215_inst_req_1 : boolean;
  signal type_cast_2215_inst_ack_1 : boolean;
  signal if_stmt_2416_branch_ack_0 : boolean;
  signal type_cast_2225_inst_req_0 : boolean;
  signal if_stmt_2379_branch_req_0 : boolean;
  signal type_cast_2225_inst_ack_0 : boolean;
  signal type_cast_2225_inst_req_1 : boolean;
  signal type_cast_2225_inst_ack_1 : boolean;
  signal addr_of_2472_final_reg_ack_0 : boolean;
  signal ptr_deref_2559_load_0_ack_0 : boolean;
  signal addr_of_2472_final_reg_req_0 : boolean;
  signal if_stmt_2416_branch_ack_1 : boolean;
  signal type_cast_2235_inst_req_0 : boolean;
  signal type_cast_2235_inst_ack_0 : boolean;
  signal type_cast_2235_inst_req_1 : boolean;
  signal type_cast_2235_inst_ack_1 : boolean;
  signal type_cast_2239_inst_req_0 : boolean;
  signal type_cast_2239_inst_ack_0 : boolean;
  signal type_cast_2239_inst_req_1 : boolean;
  signal array_obj_ref_2579_index_offset_req_0 : boolean;
  signal array_obj_ref_2579_index_offset_ack_0 : boolean;
  signal array_obj_ref_2579_index_offset_req_1 : boolean;
  signal array_obj_ref_2579_index_offset_ack_1 : boolean;
  signal addr_of_2580_final_reg_req_0 : boolean;
  signal addr_of_2580_final_reg_ack_0 : boolean;
  signal addr_of_2580_final_reg_req_1 : boolean;
  signal addr_of_2580_final_reg_ack_1 : boolean;
  signal ptr_deref_2583_store_0_req_0 : boolean;
  signal ptr_deref_2583_store_0_ack_0 : boolean;
  signal ptr_deref_2583_store_0_req_1 : boolean;
  signal ptr_deref_2583_store_0_ack_1 : boolean;
  signal type_cast_2591_inst_req_0 : boolean;
  signal type_cast_2591_inst_ack_0 : boolean;
  signal type_cast_2591_inst_req_1 : boolean;
  signal type_cast_2591_inst_ack_1 : boolean;
  signal if_stmt_2606_branch_req_0 : boolean;
  signal if_stmt_2606_branch_ack_1 : boolean;
  signal if_stmt_2606_branch_ack_0 : boolean;
  signal type_cast_2630_inst_req_0 : boolean;
  signal type_cast_2630_inst_ack_0 : boolean;
  signal type_cast_2630_inst_req_1 : boolean;
  signal type_cast_2630_inst_ack_1 : boolean;
  signal type_cast_2639_inst_req_0 : boolean;
  signal type_cast_2639_inst_ack_0 : boolean;
  signal type_cast_2639_inst_req_1 : boolean;
  signal type_cast_2639_inst_ack_1 : boolean;
  signal type_cast_2655_inst_req_0 : boolean;
  signal type_cast_2655_inst_ack_0 : boolean;
  signal type_cast_2655_inst_req_1 : boolean;
  signal type_cast_2655_inst_ack_1 : boolean;
  signal if_stmt_2662_branch_req_0 : boolean;
  signal if_stmt_2662_branch_ack_1 : boolean;
  signal if_stmt_2662_branch_ack_0 : boolean;
  signal WPIPE_Block3_complete_2692_inst_req_0 : boolean;
  signal WPIPE_Block3_complete_2692_inst_ack_0 : boolean;
  signal WPIPE_Block3_complete_2692_inst_req_1 : boolean;
  signal WPIPE_Block3_complete_2692_inst_ack_1 : boolean;
  signal phi_stmt_2329_req_0 : boolean;
  signal type_cast_2341_inst_req_0 : boolean;
  signal type_cast_2341_inst_ack_0 : boolean;
  signal type_cast_2341_inst_req_1 : boolean;
  signal type_cast_2341_inst_ack_1 : boolean;
  signal phi_stmt_2336_req_1 : boolean;
  signal type_cast_2347_inst_req_0 : boolean;
  signal type_cast_2347_inst_ack_0 : boolean;
  signal type_cast_2347_inst_req_1 : boolean;
  signal type_cast_2347_inst_ack_1 : boolean;
  signal phi_stmt_2342_req_1 : boolean;
  signal type_cast_2335_inst_req_0 : boolean;
  signal type_cast_2335_inst_ack_0 : boolean;
  signal type_cast_2335_inst_req_1 : boolean;
  signal type_cast_2335_inst_ack_1 : boolean;
  signal phi_stmt_2329_req_1 : boolean;
  signal type_cast_2339_inst_req_0 : boolean;
  signal type_cast_2339_inst_ack_0 : boolean;
  signal type_cast_2339_inst_req_1 : boolean;
  signal type_cast_2339_inst_ack_1 : boolean;
  signal phi_stmt_2336_req_0 : boolean;
  signal type_cast_2345_inst_req_0 : boolean;
  signal type_cast_2345_inst_ack_0 : boolean;
  signal type_cast_2345_inst_req_1 : boolean;
  signal type_cast_2345_inst_ack_1 : boolean;
  signal phi_stmt_2342_req_0 : boolean;
  signal phi_stmt_2329_ack_0 : boolean;
  signal phi_stmt_2336_ack_0 : boolean;
  signal phi_stmt_2342_ack_0 : boolean;
  signal phi_stmt_2669_req_1 : boolean;
  signal type_cast_2681_inst_req_0 : boolean;
  signal type_cast_2681_inst_ack_0 : boolean;
  signal type_cast_2681_inst_req_1 : boolean;
  signal type_cast_2681_inst_ack_1 : boolean;
  signal phi_stmt_2676_req_1 : boolean;
  signal type_cast_2687_inst_req_0 : boolean;
  signal type_cast_2687_inst_ack_0 : boolean;
  signal type_cast_2687_inst_req_1 : boolean;
  signal type_cast_2687_inst_ack_1 : boolean;
  signal phi_stmt_2682_req_1 : boolean;
  signal type_cast_2672_inst_req_0 : boolean;
  signal type_cast_2672_inst_ack_0 : boolean;
  signal type_cast_2672_inst_req_1 : boolean;
  signal type_cast_2672_inst_ack_1 : boolean;
  signal phi_stmt_2669_req_0 : boolean;
  signal type_cast_2679_inst_req_0 : boolean;
  signal type_cast_2679_inst_ack_0 : boolean;
  signal type_cast_2679_inst_req_1 : boolean;
  signal type_cast_2679_inst_ack_1 : boolean;
  signal phi_stmt_2676_req_0 : boolean;
  signal type_cast_2685_inst_req_0 : boolean;
  signal type_cast_2685_inst_ack_0 : boolean;
  signal type_cast_2685_inst_req_1 : boolean;
  signal type_cast_2685_inst_ack_1 : boolean;
  signal phi_stmt_2682_req_0 : boolean;
  signal phi_stmt_2669_ack_0 : boolean;
  signal phi_stmt_2676_ack_0 : boolean;
  signal phi_stmt_2682_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_D_CP_5481_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_D_CP_5481_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_D_CP_5481_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_D_CP_5481_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_D_CP_5481: Block -- control-path 
    signal zeropad3D_D_CP_5481_elements: BooleanArray(138 downto 0);
    -- 
  begin -- 
    zeropad3D_D_CP_5481_elements(0) <= zeropad3D_D_CP_5481_start;
    zeropad3D_D_CP_5481_symbol <= zeropad3D_D_CP_5481_elements(90);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2190/$entry
      -- CP-element group 0: 	 branch_block_stmt_2190/branch_block_stmt_2190__entry__
      -- CP-element group 0: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211__entry__
      -- CP-element group 0: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/$entry
      -- CP-element group 0: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_Sample/rr
      -- 
    rr_5547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(0), ack => RPIPE_Block3_starting_2192_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	138 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	99 
    -- CP-element group 1: 	100 
    -- CP-element group 1: 	102 
    -- CP-element group 1: 	103 
    -- CP-element group 1: 	105 
    -- CP-element group 1: 	106 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_2190/merge_stmt_2668__exit__
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/SplitProtocol/Update/cr
      -- 
    rr_6412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(1), ack => type_cast_2335_inst_req_0); -- 
    cr_6417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(1), ack => type_cast_2335_inst_req_1); -- 
    rr_6435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(1), ack => type_cast_2339_inst_req_0); -- 
    cr_6440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(1), ack => type_cast_2339_inst_req_1); -- 
    rr_6458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(1), ack => type_cast_2345_inst_req_0); -- 
    cr_6463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(1), ack => type_cast_2345_inst_req_1); -- 
    zeropad3D_D_CP_5481_elements(1) <= zeropad3D_D_CP_5481_elements(138);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_Update/cr
      -- 
    ra_5548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2192_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(2)); -- 
    cr_5552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(2), ack => RPIPE_Block3_starting_2192_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2192_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_Sample/rr
      -- 
    ca_5553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2192_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(3)); -- 
    rr_5561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(3), ack => RPIPE_Block3_starting_2195_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_Update/cr
      -- 
    ra_5562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2195_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(4)); -- 
    cr_5566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(4), ack => RPIPE_Block3_starting_2195_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2195_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_Sample/rr
      -- 
    ca_5567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2195_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(5)); -- 
    rr_5575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(5), ack => RPIPE_Block3_starting_2198_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_Update/cr
      -- 
    ra_5576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2198_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(6)); -- 
    cr_5580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(6), ack => RPIPE_Block3_starting_2198_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2198_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_Sample/rr
      -- 
    ca_5581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2198_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(7)); -- 
    rr_5589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(7), ack => RPIPE_Block3_starting_2201_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_Update/cr
      -- 
    ra_5590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2201_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(8)); -- 
    cr_5594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(8), ack => RPIPE_Block3_starting_2201_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2201_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_Sample/rr
      -- 
    ca_5595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2201_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(9)); -- 
    rr_5603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(9), ack => RPIPE_Block3_starting_2204_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_Update/cr
      -- 
    ra_5604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2204_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(10)); -- 
    cr_5608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(10), ack => RPIPE_Block3_starting_2204_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2204_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_Sample/rr
      -- 
    ca_5609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2204_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(11)); -- 
    rr_5617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(11), ack => RPIPE_Block3_starting_2207_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_Update/cr
      -- 
    ra_5618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2207_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(12)); -- 
    cr_5622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(12), ack => RPIPE_Block3_starting_2207_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2207_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_Sample/rr
      -- 
    ca_5623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2207_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(13)); -- 
    rr_5631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(13), ack => RPIPE_Block3_starting_2210_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_Update/cr
      -- 
    ra_5632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2210_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(14)); -- 
    cr_5636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(14), ack => RPIPE_Block3_starting_2210_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	33 
    -- CP-element group 15: 	32 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	30 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15:  members (61) 
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211__exit__
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326__entry__
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/$exit
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2193_to_assign_stmt_2211/RPIPE_Block3_starting_2210_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_Update/cr
      -- 
    ca_5637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_starting_2210_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(15)); -- 
    rr_5704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2243_inst_req_0); -- 
    cr_5751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2260_inst_req_1); -- 
    cr_5709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2243_inst_req_1); -- 
    cr_5737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2256_inst_req_1); -- 
    cr_5723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2247_inst_req_1); -- 
    rr_5718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2247_inst_req_0); -- 
    rr_5746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2260_inst_req_0); -- 
    rr_5732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2256_inst_req_0); -- 
    cr_5765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2290_inst_req_1); -- 
    rr_5760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2290_inst_req_0); -- 
    rr_5648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2215_inst_req_0); -- 
    cr_5653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2215_inst_req_1); -- 
    rr_5662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2225_inst_req_0); -- 
    cr_5667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2225_inst_req_1); -- 
    rr_5676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2235_inst_req_0); -- 
    cr_5681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2235_inst_req_1); -- 
    rr_5690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2239_inst_req_0); -- 
    cr_5695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(15), ack => type_cast_2239_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_Sample/ra
      -- 
    ra_5649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2215_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	34 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2215_Update/ca
      -- 
    ca_5654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2215_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_Sample/ra
      -- 
    ra_5663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2225_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	34 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2225_Update/ca
      -- 
    ca_5668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2225_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_Sample/ra
      -- 
    ra_5677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2235_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	34 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2235_Update/ca
      -- 
    ca_5682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2235_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_Sample/ra
      -- 
    ra_5691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2239_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2239_Update/$exit
      -- 
    ca_5696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2239_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_sample_completed_
      -- 
    ra_5705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2243_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	34 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2243_Update/ca
      -- 
    ca_5710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2243_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_sample_completed_
      -- 
    ra_5719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2247_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2247_Update/ca
      -- 
    ca_5724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2247_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_sample_completed_
      -- 
    ra_5733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2256_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2256_update_completed_
      -- 
    ca_5738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2256_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_sample_completed_
      -- 
    ra_5747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2260_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2260_update_completed_
      -- 
    ca_5752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2260_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	15 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_sample_completed_
      -- 
    ra_5761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2290_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	15 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/type_cast_2290_update_completed_
      -- 
    ca_5766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2290_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	25 
    -- CP-element group 34: 	21 
    -- CP-element group 34: 	33 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	17 
    -- CP-element group 34: 	19 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	91 
    -- CP-element group 34: 	92 
    -- CP-element group 34: 	93 
    -- CP-element group 34: 	95 
    -- CP-element group 34: 	96 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326__exit__
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody
      -- CP-element group 34: 	 branch_block_stmt_2190/assign_stmt_2216_to_assign_stmt_2326/$exit
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2329/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/SplitProtocol/Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/SplitProtocol/Update/cr
      -- 
    rr_6363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(34), ack => type_cast_2341_inst_req_0); -- 
    cr_6368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(34), ack => type_cast_2341_inst_req_1); -- 
    rr_6386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(34), ack => type_cast_2347_inst_req_0); -- 
    cr_6391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(34), ack => type_cast_2347_inst_req_1); -- 
    zeropad3D_D_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(25) & zeropad3D_D_CP_5481_elements(21) & zeropad3D_D_CP_5481_elements(33) & zeropad3D_D_CP_5481_elements(31) & zeropad3D_D_CP_5481_elements(29) & zeropad3D_D_CP_5481_elements(27) & zeropad3D_D_CP_5481_elements(23) & zeropad3D_D_CP_5481_elements(17) & zeropad3D_D_CP_5481_elements(19);
      gj_zeropad3D_D_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	113 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_Sample/$exit
      -- 
    ra_5778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2352_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(35)); -- 
    -- CP-element group 36:  branch  transition  place  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	113 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (13) 
      -- CP-element group 36: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2190/if_stmt_2379_dead_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378__exit__
      -- CP-element group 36: 	 branch_block_stmt_2190/if_stmt_2379__entry__
      -- CP-element group 36: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/$exit
      -- CP-element group 36: 	 branch_block_stmt_2190/if_stmt_2379_else_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_2190/if_stmt_2379_if_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_2190/if_stmt_2379_eval_test/branch_req
      -- CP-element group 36: 	 branch_block_stmt_2190/if_stmt_2379_eval_test/$exit
      -- CP-element group 36: 	 branch_block_stmt_2190/R_orx_xcond_2380_place
      -- CP-element group 36: 	 branch_block_stmt_2190/if_stmt_2379_eval_test/$entry
      -- 
    ca_5783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2352_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(36)); -- 
    branch_req_5791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(36), ack => if_stmt_2379_branch_req_0); -- 
    -- CP-element group 37:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	40 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (18) 
      -- CP-element group 37: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_2190/merge_stmt_2385__exit__
      -- CP-element group 37: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415__entry__
      -- CP-element group 37: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/$entry
      -- CP-element group 37: 	 branch_block_stmt_2190/if_stmt_2379_if_link/if_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_2190/if_stmt_2379_if_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_2190/whilex_xbody_lorx_xlhsx_xfalse63
      -- CP-element group 37: 	 branch_block_stmt_2190/whilex_xbody_lorx_xlhsx_xfalse63_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_2190/whilex_xbody_lorx_xlhsx_xfalse63_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_2190/merge_stmt_2385_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_2190/merge_stmt_2385_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_2190/merge_stmt_2385_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_2190/merge_stmt_2385_PhiAck/dummy
      -- 
    if_choice_transition_5796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2379_branch_ack_1, ack => zeropad3D_D_CP_5481_elements(37)); -- 
    cr_5818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(37), ack => type_cast_2389_inst_req_1); -- 
    rr_5813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(37), ack => type_cast_2389_inst_req_0); -- 
    -- CP-element group 38:  transition  place  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	114 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_2190/if_stmt_2379_else_link/else_choice_transition
      -- CP-element group 38: 	 branch_block_stmt_2190/if_stmt_2379_else_link/$exit
      -- CP-element group 38: 	 branch_block_stmt_2190/whilex_xbody_ifx_xthen
      -- CP-element group 38: 	 branch_block_stmt_2190/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_2190/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_5800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2379_branch_ack_0, ack => zeropad3D_D_CP_5481_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_sample_completed_
      -- 
    ra_5814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2389_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(39)); -- 
    -- CP-element group 40:  branch  transition  place  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	37 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (13) 
      -- CP-element group 40: 	 branch_block_stmt_2190/if_stmt_2416_eval_test/$entry
      -- CP-element group 40: 	 branch_block_stmt_2190/if_stmt_2416_eval_test/$exit
      -- CP-element group 40: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2190/if_stmt_2416_dead_link/$entry
      -- CP-element group 40: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2190/if_stmt_2416_eval_test/branch_req
      -- CP-element group 40: 	 branch_block_stmt_2190/if_stmt_2416_if_link/$entry
      -- CP-element group 40: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415__exit__
      -- CP-element group 40: 	 branch_block_stmt_2190/if_stmt_2416__entry__
      -- CP-element group 40: 	 branch_block_stmt_2190/R_orx_xcond192_2417_place
      -- CP-element group 40: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/type_cast_2389_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2190/assign_stmt_2390_to_assign_stmt_2415/$exit
      -- CP-element group 40: 	 branch_block_stmt_2190/if_stmt_2416_else_link/$entry
      -- 
    ca_5819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2389_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(40)); -- 
    branch_req_5827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(40), ack => if_stmt_2416_branch_req_0); -- 
    -- CP-element group 41:  fork  transition  place  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	57 
    -- CP-element group 41: 	58 
    -- CP-element group 41: 	60 
    -- CP-element group 41: 	62 
    -- CP-element group 41: 	64 
    -- CP-element group 41: 	66 
    -- CP-element group 41: 	68 
    -- CP-element group 41: 	70 
    -- CP-element group 41: 	72 
    -- CP-element group 41: 	75 
    -- CP-element group 41:  members (46) 
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_final_index_sum_regn_Update/req
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_final_index_sum_regn_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_complete/req
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_final_index_sum_regn_update_start
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_2190/merge_stmt_2480__exit__
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585__entry__
      -- CP-element group 41: 	 branch_block_stmt_2190/lorx_xlhsx_xfalse63_ifx_xelse
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/if_stmt_2416_if_link/if_choice_transition
      -- CP-element group 41: 	 branch_block_stmt_2190/if_stmt_2416_if_link/$exit
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_final_index_sum_regn_update_start
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_final_index_sum_regn_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_final_index_sum_regn_Update/req
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_complete/req
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_2190/lorx_xlhsx_xfalse63_ifx_xelse_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/lorx_xlhsx_xfalse63_ifx_xelse_PhiReq/$exit
      -- CP-element group 41: 	 branch_block_stmt_2190/merge_stmt_2480_PhiReqMerge
      -- CP-element group 41: 	 branch_block_stmt_2190/merge_stmt_2480_PhiAck/$entry
      -- CP-element group 41: 	 branch_block_stmt_2190/merge_stmt_2480_PhiAck/$exit
      -- CP-element group 41: 	 branch_block_stmt_2190/merge_stmt_2480_PhiAck/dummy
      -- 
    if_choice_transition_5832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2416_branch_ack_1, ack => zeropad3D_D_CP_5481_elements(41)); -- 
    req_6040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(41), ack => array_obj_ref_2554_index_offset_req_1); -- 
    req_6055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(41), ack => addr_of_2555_final_reg_req_1); -- 
    rr_5990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(41), ack => type_cast_2484_inst_req_0); -- 
    cr_6009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(41), ack => type_cast_2548_inst_req_1); -- 
    cr_5995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(41), ack => type_cast_2484_inst_req_1); -- 
    cr_6100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(41), ack => ptr_deref_2559_load_0_req_1); -- 
    cr_6119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(41), ack => type_cast_2573_inst_req_1); -- 
    req_6150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(41), ack => array_obj_ref_2579_index_offset_req_1); -- 
    req_6165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(41), ack => addr_of_2580_final_reg_req_1); -- 
    cr_6215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(41), ack => ptr_deref_2583_store_0_req_1); -- 
    -- CP-element group 42:  transition  place  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	114 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_2190/lorx_xlhsx_xfalse63_ifx_xthen
      -- CP-element group 42: 	 branch_block_stmt_2190/if_stmt_2416_else_link/else_choice_transition
      -- CP-element group 42: 	 branch_block_stmt_2190/if_stmt_2416_else_link/$exit
      -- CP-element group 42: 	 branch_block_stmt_2190/lorx_xlhsx_xfalse63_ifx_xthen_PhiReq/$entry
      -- CP-element group 42: 	 branch_block_stmt_2190/lorx_xlhsx_xfalse63_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_5836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2416_branch_ack_0, ack => zeropad3D_D_CP_5481_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	114 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_Sample/$exit
      -- 
    ra_5850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2426_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	114 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_Update/$exit
      -- 
    ca_5855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2426_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	114 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_Sample/$exit
      -- 
    ra_5864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2431_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	114 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_update_completed_
      -- 
    ca_5869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2431_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_Sample/rr
      -- CP-element group 47: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_Sample/$entry
      -- 
    rr_5877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(47), ack => type_cast_2465_inst_req_0); -- 
    zeropad3D_D_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(46) & zeropad3D_D_CP_5481_elements(44);
      gj_zeropad3D_D_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_Sample/$exit
      -- 
    ra_5878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2465_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	114 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_final_index_sum_regn_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_update_completed_
      -- 
    ca_5883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2465_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(49)); -- 
    req_5908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(49), ack => array_obj_ref_2471_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	56 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_final_index_sum_regn_Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_final_index_sum_regn_sample_complete
      -- 
    ack_5909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2471_index_offset_ack_0, ack => zeropad3D_D_CP_5481_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	114 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_request/req
      -- CP-element group 51: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_request/$entry
      -- 
    ack_5914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2471_index_offset_ack_1, ack => zeropad3D_D_CP_5481_elements(51)); -- 
    req_5923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(51), ack => addr_of_2472_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_request/ack
      -- CP-element group 52: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_request/$exit
      -- 
    ack_5924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2472_final_reg_ack_0, ack => zeropad3D_D_CP_5481_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	114 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (28) 
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/ptr_deref_2475_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/ptr_deref_2475_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/ptr_deref_2475_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/ptr_deref_2475_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/word_access_start/word_0/rr
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_base_plus_offset/$exit
      -- 
    ack_5929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2472_final_reg_ack_1, ack => zeropad3D_D_CP_5481_elements(53)); -- 
    rr_5967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(53), ack => ptr_deref_2475_store_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/word_access_start/word_0/ra
      -- CP-element group 54: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Sample/word_access_start/$exit
      -- 
    ra_5968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2475_store_0_ack_0, ack => zeropad3D_D_CP_5481_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	114 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_update_completed_
      -- 
    ca_5979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2475_store_0_ack_1, ack => zeropad3D_D_CP_5481_elements(55)); -- 
    -- CP-element group 56:  join  transition  place  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: 	50 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	115 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478__exit__
      -- CP-element group 56: 	 branch_block_stmt_2190/ifx_xthen_ifx_xend
      -- CP-element group 56: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/$exit
      -- CP-element group 56: 	 branch_block_stmt_2190/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2190/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(55) & zeropad3D_D_CP_5481_elements(50);
      gj_zeropad3D_D_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_Sample/ra
      -- 
    ra_5991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2484_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(57)); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	67 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2484_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_Sample/rr
      -- 
    ca_5996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2484_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(58)); -- 
    rr_6004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(58), ack => type_cast_2548_inst_req_0); -- 
    rr_6114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(58), ack => type_cast_2573_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_Sample/ra
      -- 
    ra_6005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2548_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	41 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (16) 
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_resized_1
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_scaled_1
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_computed_1
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_scale_1/scale_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_final_index_sum_regn_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_final_index_sum_regn_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2548_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_resize_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_resize_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_resize_1/index_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_resize_1/index_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_scale_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_scale_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_index_scale_1/scale_rename_req
      -- 
    ca_6010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2548_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(60)); -- 
    req_6035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(60), ack => array_obj_ref_2554_index_offset_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	76 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_final_index_sum_regn_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_final_index_sum_regn_sample_complete
      -- CP-element group 61: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_final_index_sum_regn_Sample/$exit
      -- 
    ack_6036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2554_index_offset_ack_0, ack => zeropad3D_D_CP_5481_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	41 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (11) 
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_request/$entry
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_final_index_sum_regn_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_final_index_sum_regn_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2554_offset_calculated
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_request/req
      -- CP-element group 62: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_sample_start_
      -- 
    ack_6041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2554_index_offset_ack_1, ack => zeropad3D_D_CP_5481_elements(62)); -- 
    req_6050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(62), ack => addr_of_2555_final_reg_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_request/$exit
      -- CP-element group 63: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_request/ack
      -- 
    ack_6051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2555_final_reg_ack_0, ack => zeropad3D_D_CP_5481_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	41 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (24) 
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_base_plus_offset/sum_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_complete/ack
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_word_addrgen/$entry
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_word_addrgen/$exit
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2555_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_base_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_word_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_root_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Sample/word_access_start/$entry
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_base_address_resized
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_base_addr_resize/$entry
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_base_addr_resize/$exit
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_base_plus_offset/sum_rename_req
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_word_addrgen/root_register_req
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_base_plus_offset/$entry
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_base_plus_offset/$exit
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Sample/word_access_start/word_0/rr
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Sample/word_access_start/word_0/$entry
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_base_addr_resize/base_resize_req
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_base_addr_resize/base_resize_ack
      -- CP-element group 64: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_word_addrgen/root_register_ack
      -- 
    ack_6056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2555_final_reg_ack_1, ack => zeropad3D_D_CP_5481_elements(64)); -- 
    rr_6089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(64), ack => ptr_deref_2559_load_0_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Sample/word_access_start/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Sample/word_access_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Sample/word_access_start/word_0/ra
      -- 
    ra_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2559_load_0_ack_0, ack => zeropad3D_D_CP_5481_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	41 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	73 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/word_access_complete/word_0/ca
      -- CP-element group 66: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/word_access_complete/word_0/$exit
      -- CP-element group 66: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/ptr_deref_2559_Merge/merge_ack
      -- CP-element group 66: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/ptr_deref_2559_Merge/$entry
      -- CP-element group 66: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/ptr_deref_2559_Merge/$exit
      -- CP-element group 66: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/ptr_deref_2559_Merge/merge_req
      -- CP-element group 66: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2559_Update/word_access_complete/$exit
      -- 
    ca_6101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2559_load_0_ack_1, ack => zeropad3D_D_CP_5481_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	58 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_Sample/ra
      -- 
    ra_6115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2573_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(67)); -- 
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	41 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/type_cast_2573_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_resized_1
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_scaled_1
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_computed_1
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_resize_1/$entry
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_resize_1/$exit
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_resize_1/index_resize_req
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_resize_1/index_resize_ack
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_scale_1/$entry
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_scale_1/$exit
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_scale_1/scale_rename_req
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_index_scale_1/scale_rename_ack
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_final_index_sum_regn_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_final_index_sum_regn_Sample/req
      -- 
    ca_6120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2573_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(68)); -- 
    req_6145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(68), ack => array_obj_ref_2579_index_offset_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	76 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_final_index_sum_regn_sample_complete
      -- CP-element group 69: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_final_index_sum_regn_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_final_index_sum_regn_Sample/ack
      -- 
    ack_6146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2579_index_offset_ack_0, ack => zeropad3D_D_CP_5481_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	41 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (11) 
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_request/$entry
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_offset_calculated
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_final_index_sum_regn_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_final_index_sum_regn_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/array_obj_ref_2579_base_plus_offset/sum_rename_ack
      -- CP-element group 70: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_request/req
      -- 
    ack_6151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2579_index_offset_ack_1, ack => zeropad3D_D_CP_5481_elements(70)); -- 
    req_6160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(70), ack => addr_of_2580_final_reg_req_0); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_request/$exit
      -- CP-element group 71: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_request/ack
      -- 
    ack_6161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2580_final_reg_ack_0, ack => zeropad3D_D_CP_5481_elements(71)); -- 
    -- CP-element group 72:  fork  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	41 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (19) 
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_complete/$exit
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/addr_of_2580_complete/ack
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_base_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_base_address_resized
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_base_addr_resize/$entry
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_base_addr_resize/$exit
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_base_addr_resize/base_resize_req
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_base_addr_resize/base_resize_ack
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_base_plus_offset/$entry
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_base_plus_offset/$exit
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_word_addrgen/$entry
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_word_addrgen/$exit
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_word_addrgen/root_register_req
      -- CP-element group 72: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_word_addrgen/root_register_ack
      -- 
    ack_6166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2580_final_reg_ack_1, ack => zeropad3D_D_CP_5481_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	66 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/ptr_deref_2583_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/ptr_deref_2583_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/ptr_deref_2583_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/ptr_deref_2583_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/word_access_start/word_0/rr
      -- 
    rr_6204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(73), ack => ptr_deref_2583_store_0_req_0); -- 
    zeropad3D_D_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(66) & zeropad3D_D_CP_5481_elements(72);
      gj_zeropad3D_D_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Sample/word_access_start/word_0/ra
      -- 
    ra_6205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2583_store_0_ack_0, ack => zeropad3D_D_CP_5481_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/ptr_deref_2583_Update/word_access_complete/word_0/ca
      -- 
    ca_6216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2583_store_0_ack_1, ack => zeropad3D_D_CP_5481_elements(75)); -- 
    -- CP-element group 76:  join  transition  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	61 
    -- CP-element group 76: 	69 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	115 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585/$exit
      -- CP-element group 76: 	 branch_block_stmt_2190/assign_stmt_2485_to_assign_stmt_2585__exit__
      -- CP-element group 76: 	 branch_block_stmt_2190/ifx_xelse_ifx_xend
      -- CP-element group 76: 	 branch_block_stmt_2190/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2190/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(61) & zeropad3D_D_CP_5481_elements(69) & zeropad3D_D_CP_5481_elements(75);
      gj_zeropad3D_D_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	115 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_Sample/ra
      -- 
    ra_6228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2591_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(77)); -- 
    -- CP-element group 78:  branch  transition  place  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	115 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (13) 
      -- CP-element group 78: 	 branch_block_stmt_2190/R_cmp147_2607_place
      -- CP-element group 78: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605__exit__
      -- CP-element group 78: 	 branch_block_stmt_2190/if_stmt_2606__entry__
      -- CP-element group 78: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/$exit
      -- CP-element group 78: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_2190/if_stmt_2606_dead_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_2190/if_stmt_2606_eval_test/$entry
      -- CP-element group 78: 	 branch_block_stmt_2190/if_stmt_2606_eval_test/$exit
      -- CP-element group 78: 	 branch_block_stmt_2190/if_stmt_2606_eval_test/branch_req
      -- CP-element group 78: 	 branch_block_stmt_2190/if_stmt_2606_if_link/$entry
      -- CP-element group 78: 	 branch_block_stmt_2190/if_stmt_2606_else_link/$entry
      -- 
    ca_6233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2591_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(78)); -- 
    branch_req_6241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(78), ack => if_stmt_2606_branch_req_0); -- 
    -- CP-element group 79:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	124 
    -- CP-element group 79: 	125 
    -- CP-element group 79: 	127 
    -- CP-element group 79: 	128 
    -- CP-element group 79: 	130 
    -- CP-element group 79: 	131 
    -- CP-element group 79:  members (40) 
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xend_ifx_xthen149
      -- CP-element group 79: 	 branch_block_stmt_2190/merge_stmt_2612__exit__
      -- CP-element group 79: 	 branch_block_stmt_2190/assign_stmt_2618__entry__
      -- CP-element group 79: 	 branch_block_stmt_2190/assign_stmt_2618__exit__
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186
      -- CP-element group 79: 	 branch_block_stmt_2190/if_stmt_2606_if_link/$exit
      -- CP-element group 79: 	 branch_block_stmt_2190/if_stmt_2606_if_link/if_choice_transition
      -- CP-element group 79: 	 branch_block_stmt_2190/assign_stmt_2618/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/assign_stmt_2618/$exit
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xend_ifx_xthen149_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xend_ifx_xthen149_PhiReq/$exit
      -- CP-element group 79: 	 branch_block_stmt_2190/merge_stmt_2612_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_2190/merge_stmt_2612_PhiAck/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/merge_stmt_2612_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_2190/merge_stmt_2612_PhiAck/dummy
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/SplitProtocol/Update/cr
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/SplitProtocol/Update/cr
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/SplitProtocol/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/SplitProtocol/Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/SplitProtocol/Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/SplitProtocol/Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2606_branch_ack_1, ack => zeropad3D_D_CP_5481_elements(79)); -- 
    rr_6618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(79), ack => type_cast_2672_inst_req_0); -- 
    cr_6623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(79), ack => type_cast_2672_inst_req_1); -- 
    rr_6641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(79), ack => type_cast_2679_inst_req_0); -- 
    cr_6646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(79), ack => type_cast_2679_inst_req_1); -- 
    rr_6664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(79), ack => type_cast_2685_inst_req_0); -- 
    cr_6669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(79), ack => type_cast_2685_inst_req_1); -- 
    -- CP-element group 80:  fork  transition  place  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80: 	84 
    -- CP-element group 80: 	86 
    -- CP-element group 80:  members (24) 
      -- CP-element group 80: 	 branch_block_stmt_2190/ifx_xend_ifx_xelse154
      -- CP-element group 80: 	 branch_block_stmt_2190/merge_stmt_2620__exit__
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661__entry__
      -- CP-element group 80: 	 branch_block_stmt_2190/if_stmt_2606_else_link/$exit
      -- CP-element group 80: 	 branch_block_stmt_2190/if_stmt_2606_else_link/else_choice_transition
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/$entry
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_update_start_
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_update_start_
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_update_start_
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_2190/ifx_xend_ifx_xelse154_PhiReq/$entry
      -- CP-element group 80: 	 branch_block_stmt_2190/ifx_xend_ifx_xelse154_PhiReq/$exit
      -- CP-element group 80: 	 branch_block_stmt_2190/merge_stmt_2620_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_2190/merge_stmt_2620_PhiAck/$entry
      -- CP-element group 80: 	 branch_block_stmt_2190/merge_stmt_2620_PhiAck/$exit
      -- CP-element group 80: 	 branch_block_stmt_2190/merge_stmt_2620_PhiAck/dummy
      -- 
    else_choice_transition_6250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2606_branch_ack_0, ack => zeropad3D_D_CP_5481_elements(80)); -- 
    rr_6266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(80), ack => type_cast_2630_inst_req_0); -- 
    cr_6271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(80), ack => type_cast_2630_inst_req_1); -- 
    cr_6285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(80), ack => type_cast_2639_inst_req_1); -- 
    cr_6299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(80), ack => type_cast_2655_inst_req_1); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_Sample/ra
      -- 
    ra_6267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2630_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2630_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_Sample/rr
      -- 
    ca_6272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2630_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(82)); -- 
    rr_6280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(82), ack => type_cast_2639_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_Sample/ra
      -- 
    ra_6281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2639_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2639_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_Sample/rr
      -- 
    ca_6286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2639_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(84)); -- 
    rr_6294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(84), ack => type_cast_2655_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_Sample/ra
      -- 
    ra_6295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2655_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(85)); -- 
    -- CP-element group 86:  branch  transition  place  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	80 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (13) 
      -- CP-element group 86: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661__exit__
      -- CP-element group 86: 	 branch_block_stmt_2190/if_stmt_2662__entry__
      -- CP-element group 86: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/$exit
      -- CP-element group 86: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2190/assign_stmt_2626_to_assign_stmt_2661/type_cast_2655_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_2190/if_stmt_2662_dead_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2190/if_stmt_2662_eval_test/$entry
      -- CP-element group 86: 	 branch_block_stmt_2190/if_stmt_2662_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_2190/if_stmt_2662_eval_test/branch_req
      -- CP-element group 86: 	 branch_block_stmt_2190/R_cmp178_2663_place
      -- CP-element group 86: 	 branch_block_stmt_2190/if_stmt_2662_if_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2190/if_stmt_2662_else_link/$entry
      -- 
    ca_6300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2655_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(86)); -- 
    branch_req_6308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(86), ack => if_stmt_2662_branch_req_0); -- 
    -- CP-element group 87:  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (15) 
      -- CP-element group 87: 	 branch_block_stmt_2190/merge_stmt_2690__exit__
      -- CP-element group 87: 	 branch_block_stmt_2190/assign_stmt_2695__entry__
      -- CP-element group 87: 	 branch_block_stmt_2190/if_stmt_2662_if_link/$exit
      -- CP-element group 87: 	 branch_block_stmt_2190/if_stmt_2662_if_link/if_choice_transition
      -- CP-element group 87: 	 branch_block_stmt_2190/ifx_xelse154_whilex_xend
      -- CP-element group 87: 	 branch_block_stmt_2190/assign_stmt_2695/$entry
      -- CP-element group 87: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_Sample/req
      -- CP-element group 87: 	 branch_block_stmt_2190/ifx_xelse154_whilex_xend_PhiReq/$entry
      -- CP-element group 87: 	 branch_block_stmt_2190/ifx_xelse154_whilex_xend_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_2190/merge_stmt_2690_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_2190/merge_stmt_2690_PhiAck/$entry
      -- CP-element group 87: 	 branch_block_stmt_2190/merge_stmt_2690_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_2190/merge_stmt_2690_PhiAck/dummy
      -- 
    if_choice_transition_6313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2662_branch_ack_1, ack => zeropad3D_D_CP_5481_elements(87)); -- 
    req_6330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(87), ack => WPIPE_Block3_complete_2692_inst_req_0); -- 
    -- CP-element group 88:  fork  transition  place  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	116 
    -- CP-element group 88: 	117 
    -- CP-element group 88: 	118 
    -- CP-element group 88: 	120 
    -- CP-element group 88: 	121 
    -- CP-element group 88:  members (22) 
      -- CP-element group 88: 	 branch_block_stmt_2190/if_stmt_2662_else_link/$exit
      -- CP-element group 88: 	 branch_block_stmt_2190/if_stmt_2662_else_link/else_choice_transition
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2669/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/SplitProtocol/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/SplitProtocol/Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/SplitProtocol/Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/SplitProtocol/Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/SplitProtocol/Update/cr
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/SplitProtocol/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/SplitProtocol/Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/SplitProtocol/Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/SplitProtocol/Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2662_branch_ack_0, ack => zeropad3D_D_CP_5481_elements(88)); -- 
    rr_6569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(88), ack => type_cast_2681_inst_req_0); -- 
    cr_6574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(88), ack => type_cast_2681_inst_req_1); -- 
    rr_6592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(88), ack => type_cast_2687_inst_req_0); -- 
    cr_6597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(88), ack => type_cast_2687_inst_req_1); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_update_start_
      -- CP-element group 89: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_Sample/ack
      -- CP-element group 89: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_Update/req
      -- 
    ack_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_complete_2692_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(89)); -- 
    req_6335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(89), ack => WPIPE_Block3_complete_2692_inst_req_1); -- 
    -- CP-element group 90:  transition  place  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (16) 
      -- CP-element group 90: 	 $exit
      -- CP-element group 90: 	 branch_block_stmt_2190/$exit
      -- CP-element group 90: 	 branch_block_stmt_2190/branch_block_stmt_2190__exit__
      -- CP-element group 90: 	 branch_block_stmt_2190/assign_stmt_2695__exit__
      -- CP-element group 90: 	 branch_block_stmt_2190/return__
      -- CP-element group 90: 	 branch_block_stmt_2190/merge_stmt_2697__exit__
      -- CP-element group 90: 	 branch_block_stmt_2190/assign_stmt_2695/$exit
      -- CP-element group 90: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2190/assign_stmt_2695/WPIPE_Block3_complete_2692_Update/ack
      -- CP-element group 90: 	 branch_block_stmt_2190/return___PhiReq/$entry
      -- CP-element group 90: 	 branch_block_stmt_2190/return___PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_2190/merge_stmt_2697_PhiReqMerge
      -- CP-element group 90: 	 branch_block_stmt_2190/merge_stmt_2697_PhiAck/$entry
      -- CP-element group 90: 	 branch_block_stmt_2190/merge_stmt_2697_PhiAck/$exit
      -- CP-element group 90: 	 branch_block_stmt_2190/merge_stmt_2697_PhiAck/dummy
      -- 
    ack_6336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_complete_2692_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(90)); -- 
    -- CP-element group 91:  transition  output  delay-element  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	34 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2329/$exit
      -- CP-element group 91: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2333_konst_delay_trans
      -- CP-element group 91: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_req
      -- 
    phi_stmt_2329_req_6347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2329_req_6347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(91), ack => phi_stmt_2329_req_0); -- 
    -- Element group zeropad3D_D_CP_5481_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => zeropad3D_D_CP_5481_elements(34), ack => zeropad3D_D_CP_5481_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	34 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/SplitProtocol/Sample/ra
      -- 
    ra_6364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	34 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/SplitProtocol/Update/ca
      -- 
    ca_6369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/$exit
      -- CP-element group 94: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/$exit
      -- CP-element group 94: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2341/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_req
      -- 
    phi_stmt_2336_req_6370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2336_req_6370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(94), ack => phi_stmt_2336_req_1); -- 
    zeropad3D_D_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(92) & zeropad3D_D_CP_5481_elements(93);
      gj_zeropad3D_D_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	34 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/SplitProtocol/Sample/ra
      -- 
    ra_6387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	34 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/SplitProtocol/Update/ca
      -- 
    ca_6392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/$exit
      -- CP-element group 97: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/$exit
      -- CP-element group 97: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2347/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_req
      -- 
    phi_stmt_2342_req_6393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2342_req_6393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(97), ack => phi_stmt_2342_req_1); -- 
    zeropad3D_D_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(95) & zeropad3D_D_CP_5481_elements(96);
      gj_zeropad3D_D_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	109 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2190/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_D_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(91) & zeropad3D_D_CP_5481_elements(94) & zeropad3D_D_CP_5481_elements(97);
      gj_zeropad3D_D_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	1 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/SplitProtocol/Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/SplitProtocol/Sample/ra
      -- 
    ra_6413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2335_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	1 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/SplitProtocol/Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/SplitProtocol/Update/ca
      -- 
    ca_6418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2335_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/$exit
      -- CP-element group 101: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/$exit
      -- CP-element group 101: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_sources/type_cast_2335/SplitProtocol/$exit
      -- CP-element group 101: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2329/phi_stmt_2329_req
      -- 
    phi_stmt_2329_req_6419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2329_req_6419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(101), ack => phi_stmt_2329_req_1); -- 
    zeropad3D_D_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(99) & zeropad3D_D_CP_5481_elements(100);
      gj_zeropad3D_D_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	1 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/SplitProtocol/Sample/ra
      -- 
    ra_6436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2339_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	1 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/SplitProtocol/Update/ca
      -- 
    ca_6441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2339_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/$exit
      -- CP-element group 104: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/$exit
      -- CP-element group 104: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_sources/type_cast_2339/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2336/phi_stmt_2336_req
      -- 
    phi_stmt_2336_req_6442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2336_req_6442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(104), ack => phi_stmt_2336_req_0); -- 
    zeropad3D_D_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(102) & zeropad3D_D_CP_5481_elements(103);
      gj_zeropad3D_D_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	1 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/SplitProtocol/Sample/ra
      -- 
    ra_6459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2345_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	1 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/SplitProtocol/Update/ca
      -- 
    ca_6464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2345_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/$exit
      -- CP-element group 107: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/$exit
      -- CP-element group 107: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2345/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_req
      -- 
    phi_stmt_2342_req_6465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2342_req_6465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(107), ack => phi_stmt_2342_req_0); -- 
    zeropad3D_D_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(105) & zeropad3D_D_CP_5481_elements(106);
      gj_zeropad3D_D_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2190/ifx_xend186_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(101) & zeropad3D_D_CP_5481_elements(104) & zeropad3D_D_CP_5481_elements(107);
      gj_zeropad3D_D_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  merge  fork  transition  place  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	98 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	112 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2190/merge_stmt_2328_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_2190/merge_stmt_2328_PhiAck/$entry
      -- 
    zeropad3D_D_CP_5481_elements(109) <= OrReduce(zeropad3D_D_CP_5481_elements(98) & zeropad3D_D_CP_5481_elements(108));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_2190/merge_stmt_2328_PhiAck/phi_stmt_2329_ack
      -- 
    phi_stmt_2329_ack_6470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2329_ack_0, ack => zeropad3D_D_CP_5481_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_2190/merge_stmt_2328_PhiAck/phi_stmt_2336_ack
      -- 
    phi_stmt_2336_ack_6471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2336_ack_0, ack => zeropad3D_D_CP_5481_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	109 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2190/merge_stmt_2328_PhiAck/phi_stmt_2342_ack
      -- 
    phi_stmt_2342_ack_6472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2342_ack_0, ack => zeropad3D_D_CP_5481_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  place  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	35 
    -- CP-element group 113: 	36 
    -- CP-element group 113:  members (10) 
      -- CP-element group 113: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_update_start_
      -- CP-element group 113: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_Update/cr
      -- CP-element group 113: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/type_cast_2352_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_2190/merge_stmt_2328__exit__
      -- CP-element group 113: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378__entry__
      -- CP-element group 113: 	 branch_block_stmt_2190/assign_stmt_2353_to_assign_stmt_2378/$entry
      -- CP-element group 113: 	 branch_block_stmt_2190/merge_stmt_2328_PhiAck/$exit
      -- 
    cr_5782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(113), ack => type_cast_2352_inst_req_1); -- 
    rr_5777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(113), ack => type_cast_2352_inst_req_0); -- 
    zeropad3D_D_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(110) & zeropad3D_D_CP_5481_elements(111) & zeropad3D_D_CP_5481_elements(112);
      gj_zeropad3D_D_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  merge  fork  transition  place  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	38 
    -- CP-element group 114: 	42 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	45 
    -- CP-element group 114: 	46 
    -- CP-element group 114: 	55 
    -- CP-element group 114: 	49 
    -- CP-element group 114: 	51 
    -- CP-element group 114: 	53 
    -- CP-element group 114: 	44 
    -- CP-element group 114: 	43 
    -- CP-element group 114:  members (33) 
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Update/word_access_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Update/word_access_complete/word_0/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Update/word_access_complete/word_0/cr
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_complete/req
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_final_index_sum_regn_Update/req
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_final_index_sum_regn_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/merge_stmt_2422__exit__
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478__entry__
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/array_obj_ref_2471_final_index_sum_regn_update_start
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2431_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/ptr_deref_2475_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2426_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/addr_of_2472_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/assign_stmt_2427_to_assign_stmt_2478/type_cast_2465_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2190/merge_stmt_2422_PhiReqMerge
      -- CP-element group 114: 	 branch_block_stmt_2190/merge_stmt_2422_PhiAck/$entry
      -- CP-element group 114: 	 branch_block_stmt_2190/merge_stmt_2422_PhiAck/$exit
      -- CP-element group 114: 	 branch_block_stmt_2190/merge_stmt_2422_PhiAck/dummy
      -- 
    cr_5978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(114), ack => ptr_deref_2475_store_0_req_1); -- 
    cr_5868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(114), ack => type_cast_2431_inst_req_1); -- 
    req_5928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(114), ack => addr_of_2472_final_reg_req_1); -- 
    req_5913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(114), ack => array_obj_ref_2471_index_offset_req_1); -- 
    rr_5863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(114), ack => type_cast_2431_inst_req_0); -- 
    cr_5882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(114), ack => type_cast_2465_inst_req_1); -- 
    cr_5854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(114), ack => type_cast_2426_inst_req_1); -- 
    rr_5849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(114), ack => type_cast_2426_inst_req_0); -- 
    zeropad3D_D_CP_5481_elements(114) <= OrReduce(zeropad3D_D_CP_5481_elements(38) & zeropad3D_D_CP_5481_elements(42));
    -- CP-element group 115:  merge  fork  transition  place  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	56 
    -- CP-element group 115: 	76 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	77 
    -- CP-element group 115: 	78 
    -- CP-element group 115:  members (13) 
      -- CP-element group 115: 	 branch_block_stmt_2190/merge_stmt_2587__exit__
      -- CP-element group 115: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605__entry__
      -- CP-element group 115: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/$entry
      -- CP-element group 115: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_update_start_
      -- CP-element group 115: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_2190/assign_stmt_2592_to_assign_stmt_2605/type_cast_2591_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_2190/merge_stmt_2587_PhiReqMerge
      -- CP-element group 115: 	 branch_block_stmt_2190/merge_stmt_2587_PhiAck/$entry
      -- CP-element group 115: 	 branch_block_stmt_2190/merge_stmt_2587_PhiAck/$exit
      -- CP-element group 115: 	 branch_block_stmt_2190/merge_stmt_2587_PhiAck/dummy
      -- 
    rr_6227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(115), ack => type_cast_2591_inst_req_0); -- 
    cr_6232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(115), ack => type_cast_2591_inst_req_1); -- 
    zeropad3D_D_CP_5481_elements(115) <= OrReduce(zeropad3D_D_CP_5481_elements(56) & zeropad3D_D_CP_5481_elements(76));
    -- CP-element group 116:  transition  output  delay-element  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	88 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	123 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2669/$exit
      -- CP-element group 116: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2675_konst_delay_trans
      -- CP-element group 116: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_req
      -- 
    phi_stmt_2669_req_6553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2669_req_6553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(116), ack => phi_stmt_2669_req_1); -- 
    -- Element group zeropad3D_D_CP_5481_elements(116) is a control-delay.
    cp_element_116_delay: control_delay_element  generic map(name => " 116_delay", delay_value => 1)  port map(req => zeropad3D_D_CP_5481_elements(88), ack => zeropad3D_D_CP_5481_elements(116), clk => clk, reset =>reset);
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	88 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/SplitProtocol/Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/SplitProtocol/Sample/ra
      -- 
    ra_6570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2681_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	88 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/SplitProtocol/Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/SplitProtocol/Update/ca
      -- 
    ca_6575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2681_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/$exit
      -- CP-element group 119: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/$exit
      -- CP-element group 119: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2681/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_req
      -- 
    phi_stmt_2676_req_6576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2676_req_6576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(119), ack => phi_stmt_2676_req_1); -- 
    zeropad3D_D_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(117) & zeropad3D_D_CP_5481_elements(118);
      gj_zeropad3D_D_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	88 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/SplitProtocol/Sample/ra
      -- 
    ra_6593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2687_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	88 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/SplitProtocol/Update/ca
      -- 
    ca_6598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2687_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/$exit
      -- CP-element group 122: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/$exit
      -- CP-element group 122: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2687/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_req
      -- 
    phi_stmt_2682_req_6599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2682_req_6599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(122), ack => phi_stmt_2682_req_1); -- 
    zeropad3D_D_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(120) & zeropad3D_D_CP_5481_elements(121);
      gj_zeropad3D_D_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	116 
    -- CP-element group 123: 	119 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	134 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2190/ifx_xelse154_ifx_xend186_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(116) & zeropad3D_D_CP_5481_elements(119) & zeropad3D_D_CP_5481_elements(122);
      gj_zeropad3D_D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	79 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/SplitProtocol/Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/SplitProtocol/Sample/ra
      -- 
    ra_6619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2672_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	79 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/SplitProtocol/Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/SplitProtocol/Update/ca
      -- 
    ca_6624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2672_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	133 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/$exit
      -- CP-element group 126: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/$exit
      -- CP-element group 126: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/$exit
      -- CP-element group 126: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_sources/type_cast_2672/SplitProtocol/$exit
      -- CP-element group 126: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2669/phi_stmt_2669_req
      -- 
    phi_stmt_2669_req_6625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2669_req_6625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(126), ack => phi_stmt_2669_req_0); -- 
    zeropad3D_D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(124) & zeropad3D_D_CP_5481_elements(125);
      gj_zeropad3D_D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	79 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/SplitProtocol/Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/SplitProtocol/Sample/ra
      -- 
    ra_6642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2679_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	79 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/SplitProtocol/Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/SplitProtocol/Update/ca
      -- 
    ca_6647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2679_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	133 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/$exit
      -- CP-element group 129: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/$exit
      -- CP-element group 129: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/$exit
      -- CP-element group 129: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_sources/type_cast_2679/SplitProtocol/$exit
      -- CP-element group 129: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2676/phi_stmt_2676_req
      -- 
    phi_stmt_2676_req_6648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2676_req_6648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(129), ack => phi_stmt_2676_req_0); -- 
    zeropad3D_D_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(127) & zeropad3D_D_CP_5481_elements(128);
      gj_zeropad3D_D_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	79 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/SplitProtocol/Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/SplitProtocol/Sample/ra
      -- 
    ra_6665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2685_inst_ack_0, ack => zeropad3D_D_CP_5481_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	79 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/SplitProtocol/Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/SplitProtocol/Update/ca
      -- 
    ca_6670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2685_inst_ack_1, ack => zeropad3D_D_CP_5481_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/$exit
      -- CP-element group 132: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/$exit
      -- CP-element group 132: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/$exit
      -- CP-element group 132: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_sources/type_cast_2685/SplitProtocol/$exit
      -- CP-element group 132: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/phi_stmt_2682/phi_stmt_2682_req
      -- 
    phi_stmt_2682_req_6671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2682_req_6671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_D_CP_5481_elements(132), ack => phi_stmt_2682_req_0); -- 
    zeropad3D_D_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(130) & zeropad3D_D_CP_5481_elements(131);
      gj_zeropad3D_D_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	126 
    -- CP-element group 133: 	129 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_2190/ifx_xthen149_ifx_xend186_PhiReq/$exit
      -- 
    zeropad3D_D_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(126) & zeropad3D_D_CP_5481_elements(129) & zeropad3D_D_CP_5481_elements(132);
      gj_zeropad3D_D_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  merge  fork  transition  place  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	123 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	136 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_2190/merge_stmt_2668_PhiReqMerge
      -- CP-element group 134: 	 branch_block_stmt_2190/merge_stmt_2668_PhiAck/$entry
      -- 
    zeropad3D_D_CP_5481_elements(134) <= OrReduce(zeropad3D_D_CP_5481_elements(123) & zeropad3D_D_CP_5481_elements(133));
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	138 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_2190/merge_stmt_2668_PhiAck/phi_stmt_2669_ack
      -- 
    phi_stmt_2669_ack_6676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2669_ack_0, ack => zeropad3D_D_CP_5481_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_2190/merge_stmt_2668_PhiAck/phi_stmt_2676_ack
      -- 
    phi_stmt_2676_ack_6677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2676_ack_0, ack => zeropad3D_D_CP_5481_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_2190/merge_stmt_2668_PhiAck/phi_stmt_2682_ack
      -- 
    phi_stmt_2682_ack_6678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2682_ack_0, ack => zeropad3D_D_CP_5481_elements(137)); -- 
    -- CP-element group 138:  join  transition  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: 	136 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	1 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_2190/merge_stmt_2668_PhiAck/$exit
      -- 
    zeropad3D_D_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_D_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_D_CP_5481_elements(135) & zeropad3D_D_CP_5481_elements(136) & zeropad3D_D_CP_5481_elements(137);
      gj_zeropad3D_D_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_D_CP_5481_elements(138), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2274_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2324_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2459_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2542_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2567_wire : std_logic_vector(31 downto 0);
    signal R_idxprom134_2553_resized : std_logic_vector(13 downto 0);
    signal R_idxprom134_2553_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom139_2578_resized : std_logic_vector(13 downto 0);
    signal R_idxprom139_2578_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2470_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2470_scaled : std_logic_vector(13 downto 0);
    signal add106_2510 : std_logic_vector(31 downto 0);
    signal add115_2515 : std_logic_vector(31 downto 0);
    signal add125_2530 : std_logic_vector(31 downto 0);
    signal add131_2535 : std_logic_vector(31 downto 0);
    signal add144_2598 : std_logic_vector(31 downto 0);
    signal add152_2618 : std_logic_vector(15 downto 0);
    signal add162_2287 : std_logic_vector(31 downto 0);
    signal add177_2296 : std_logic_vector(31 downto 0);
    signal add77_2306 : std_logic_vector(31 downto 0);
    signal add88_2447 : std_logic_vector(31 downto 0);
    signal add94_2452 : std_logic_vector(31 downto 0);
    signal add_2301 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2471_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2471_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2471_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2471_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2471_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2471_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2554_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2554_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2554_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2554_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2554_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2554_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2579_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2579_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2579_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2579_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2579_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2579_root_address : std_logic_vector(13 downto 0);
    signal arrayidx135_2556 : std_logic_vector(31 downto 0);
    signal arrayidx140_2581 : std_logic_vector(31 downto 0);
    signal arrayidx_2473 : std_logic_vector(31 downto 0);
    signal call1_2196 : std_logic_vector(7 downto 0);
    signal call2_2199 : std_logic_vector(7 downto 0);
    signal call3_2202 : std_logic_vector(7 downto 0);
    signal call4_2205 : std_logic_vector(7 downto 0);
    signal call5_2208 : std_logic_vector(7 downto 0);
    signal call6_2211 : std_logic_vector(7 downto 0);
    signal call_2193 : std_logic_vector(7 downto 0);
    signal cmp147_2605 : std_logic_vector(0 downto 0);
    signal cmp163_2636 : std_logic_vector(0 downto 0);
    signal cmp178_2661 : std_logic_vector(0 downto 0);
    signal cmp61_2373 : std_logic_vector(0 downto 0);
    signal cmp68_2397 : std_logic_vector(0 downto 0);
    signal cmp68x_xnot_2403 : std_logic_vector(0 downto 0);
    signal cmp78_2410 : std_logic_vector(0 downto 0);
    signal cmp_2360 : std_logic_vector(0 downto 0);
    signal cmpx_xnot_2366 : std_logic_vector(0 downto 0);
    signal conv108_2326 : std_logic_vector(31 downto 0);
    signal conv10_2226 : std_logic_vector(15 downto 0);
    signal conv143_2592 : std_logic_vector(31 downto 0);
    signal conv157_2631 : std_logic_vector(31 downto 0);
    signal conv171_2656 : std_logic_vector(31 downto 0);
    signal conv173_2291 : std_logic_vector(31 downto 0);
    signal conv36_2236 : std_logic_vector(31 downto 0);
    signal conv38_2240 : std_logic_vector(31 downto 0);
    signal conv42_2244 : std_logic_vector(31 downto 0);
    signal conv44_2248 : std_logic_vector(31 downto 0);
    signal conv51_2353 : std_logic_vector(31 downto 0);
    signal conv53_2257 : std_logic_vector(31 downto 0);
    signal conv65_2390 : std_logic_vector(31 downto 0);
    signal conv82_2427 : std_logic_vector(31 downto 0);
    signal conv84_2261 : std_logic_vector(31 downto 0);
    signal conv86_2432 : std_logic_vector(31 downto 0);
    signal conv90_2276 : std_logic_vector(31 downto 0);
    signal conv98_2485 : std_logic_vector(31 downto 0);
    signal conv_2216 : std_logic_vector(15 downto 0);
    signal div11_2232 : std_logic_vector(15 downto 0);
    signal div_2222 : std_logic_vector(15 downto 0);
    signal idxprom134_2549 : std_logic_vector(63 downto 0);
    signal idxprom139_2574 : std_logic_vector(63 downto 0);
    signal idxprom_2466 : std_logic_vector(63 downto 0);
    signal inc168_2640 : std_logic_vector(15 downto 0);
    signal inc168x_xix_x2_2645 : std_logic_vector(15 downto 0);
    signal inc_2626 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_2676 : std_logic_vector(15 downto 0);
    signal ix_x2_2336 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_2682 : std_logic_vector(15 downto 0);
    signal jx_x1_2342 : std_logic_vector(15 downto 0);
    signal jx_x2_2651 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_2669 : std_logic_vector(15 downto 0);
    signal kx_x1_2329 : std_logic_vector(15 downto 0);
    signal mul105_2495 : std_logic_vector(31 downto 0);
    signal mul114_2505 : std_logic_vector(31 downto 0);
    signal mul124_2520 : std_logic_vector(31 downto 0);
    signal mul130_2525 : std_logic_vector(31 downto 0);
    signal mul45_2253 : std_logic_vector(31 downto 0);
    signal mul87_2437 : std_logic_vector(31 downto 0);
    signal mul93_2442 : std_logic_vector(31 downto 0);
    signal mul_2312 : std_logic_vector(31 downto 0);
    signal orx_xcond192_2415 : std_logic_vector(0 downto 0);
    signal orx_xcond_2378 : std_logic_vector(0 downto 0);
    signal ptr_deref_2475_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2475_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2475_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2475_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2475_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2475_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2559_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2559_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2559_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2559_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2559_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2583_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2583_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2583_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2583_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2583_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2583_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext191_2267 : std_logic_vector(31 downto 0);
    signal sext_2317 : std_logic_vector(31 downto 0);
    signal shl_2282 : std_logic_vector(31 downto 0);
    signal shr133_2544 : std_logic_vector(31 downto 0);
    signal shr138_2569 : std_logic_vector(31 downto 0);
    signal shr_2461 : std_logic_vector(31 downto 0);
    signal sub113_2500 : std_logic_vector(31 downto 0);
    signal sub_2490 : std_logic_vector(31 downto 0);
    signal tmp136_2560 : std_logic_vector(63 downto 0);
    signal type_cast_2220_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2230_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2265_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2270_wire : std_logic_vector(31 downto 0);
    signal type_cast_2273_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2280_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2310_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2320_wire : std_logic_vector(31 downto 0);
    signal type_cast_2323_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2333_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2335_wire : std_logic_vector(15 downto 0);
    signal type_cast_2339_wire : std_logic_vector(15 downto 0);
    signal type_cast_2341_wire : std_logic_vector(15 downto 0);
    signal type_cast_2345_wire : std_logic_vector(15 downto 0);
    signal type_cast_2347_wire : std_logic_vector(15 downto 0);
    signal type_cast_2351_wire : std_logic_vector(31 downto 0);
    signal type_cast_2356_wire : std_logic_vector(31 downto 0);
    signal type_cast_2358_wire : std_logic_vector(31 downto 0);
    signal type_cast_2364_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2369_wire : std_logic_vector(31 downto 0);
    signal type_cast_2371_wire : std_logic_vector(31 downto 0);
    signal type_cast_2388_wire : std_logic_vector(31 downto 0);
    signal type_cast_2393_wire : std_logic_vector(31 downto 0);
    signal type_cast_2395_wire : std_logic_vector(31 downto 0);
    signal type_cast_2401_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2406_wire : std_logic_vector(31 downto 0);
    signal type_cast_2408_wire : std_logic_vector(31 downto 0);
    signal type_cast_2425_wire : std_logic_vector(31 downto 0);
    signal type_cast_2430_wire : std_logic_vector(31 downto 0);
    signal type_cast_2455_wire : std_logic_vector(31 downto 0);
    signal type_cast_2458_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2464_wire : std_logic_vector(63 downto 0);
    signal type_cast_2477_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2483_wire : std_logic_vector(31 downto 0);
    signal type_cast_2538_wire : std_logic_vector(31 downto 0);
    signal type_cast_2541_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2547_wire : std_logic_vector(63 downto 0);
    signal type_cast_2563_wire : std_logic_vector(31 downto 0);
    signal type_cast_2566_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2572_wire : std_logic_vector(63 downto 0);
    signal type_cast_2590_wire : std_logic_vector(31 downto 0);
    signal type_cast_2596_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2601_wire : std_logic_vector(31 downto 0);
    signal type_cast_2603_wire : std_logic_vector(31 downto 0);
    signal type_cast_2616_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2624_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2629_wire : std_logic_vector(31 downto 0);
    signal type_cast_2654_wire : std_logic_vector(31 downto 0);
    signal type_cast_2672_wire : std_logic_vector(15 downto 0);
    signal type_cast_2675_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2679_wire : std_logic_vector(15 downto 0);
    signal type_cast_2681_wire : std_logic_vector(15 downto 0);
    signal type_cast_2685_wire : std_logic_vector(15 downto 0);
    signal type_cast_2687_wire : std_logic_vector(15 downto 0);
    signal type_cast_2694_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_2471_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2471_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2471_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2471_resized_base_address <= "00000000000000";
    array_obj_ref_2554_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2554_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2554_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2554_resized_base_address <= "00000000000000";
    array_obj_ref_2579_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2579_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2579_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2579_resized_base_address <= "00000000000000";
    ptr_deref_2475_word_offset_0 <= "00000000000000";
    ptr_deref_2559_word_offset_0 <= "00000000000000";
    ptr_deref_2583_word_offset_0 <= "00000000000000";
    type_cast_2220_wire_constant <= "0000000000000001";
    type_cast_2230_wire_constant <= "0000000000000001";
    type_cast_2265_wire_constant <= "00000000000000000000000000010000";
    type_cast_2273_wire_constant <= "00000000000000000000000000010000";
    type_cast_2280_wire_constant <= "00000000000000000000000000000001";
    type_cast_2310_wire_constant <= "00000000000000000000000000010000";
    type_cast_2323_wire_constant <= "00000000000000000000000000010000";
    type_cast_2333_wire_constant <= "0000000000000000";
    type_cast_2364_wire_constant <= "1";
    type_cast_2401_wire_constant <= "1";
    type_cast_2458_wire_constant <= "00000000000000000000000000000010";
    type_cast_2477_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2541_wire_constant <= "00000000000000000000000000000010";
    type_cast_2566_wire_constant <= "00000000000000000000000000000010";
    type_cast_2596_wire_constant <= "00000000000000000000000000000100";
    type_cast_2616_wire_constant <= "0000000000000100";
    type_cast_2624_wire_constant <= "0000000000000001";
    type_cast_2675_wire_constant <= "0000000000000000";
    type_cast_2694_wire_constant <= "00000001";
    phi_stmt_2329: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2333_wire_constant & type_cast_2335_wire;
      req <= phi_stmt_2329_req_0 & phi_stmt_2329_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2329",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2329_ack_0,
          idata => idata,
          odata => kx_x1_2329,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2329
    phi_stmt_2336: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2339_wire & type_cast_2341_wire;
      req <= phi_stmt_2336_req_0 & phi_stmt_2336_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2336",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2336_ack_0,
          idata => idata,
          odata => ix_x2_2336,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2336
    phi_stmt_2342: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2345_wire & type_cast_2347_wire;
      req <= phi_stmt_2342_req_0 & phi_stmt_2342_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2342",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2342_ack_0,
          idata => idata,
          odata => jx_x1_2342,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2342
    phi_stmt_2669: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2672_wire & type_cast_2675_wire_constant;
      req <= phi_stmt_2669_req_0 & phi_stmt_2669_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2669",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2669_ack_0,
          idata => idata,
          odata => kx_x0x_xph_2669,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2669
    phi_stmt_2676: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2679_wire & type_cast_2681_wire;
      req <= phi_stmt_2676_req_0 & phi_stmt_2676_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2676",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2676_ack_0,
          idata => idata,
          odata => ix_x1x_xph_2676,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2676
    phi_stmt_2682: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2685_wire & type_cast_2687_wire;
      req <= phi_stmt_2682_req_0 & phi_stmt_2682_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2682",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2682_ack_0,
          idata => idata,
          odata => jx_x0x_xph_2682,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2682
    -- flow-through select operator MUX_2650_inst
    jx_x2_2651 <= div_2222 when (cmp163_2636(0) /=  '0') else inc_2626;
    addr_of_2472_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2472_final_reg_req_0;
      addr_of_2472_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2472_final_reg_req_1;
      addr_of_2472_final_reg_ack_1<= rack(0);
      addr_of_2472_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2472_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2471_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2555_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2555_final_reg_req_0;
      addr_of_2555_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2555_final_reg_req_1;
      addr_of_2555_final_reg_ack_1<= rack(0);
      addr_of_2555_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2555_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2554_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx135_2556,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2580_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2580_final_reg_req_0;
      addr_of_2580_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2580_final_reg_req_1;
      addr_of_2580_final_reg_ack_1<= rack(0);
      addr_of_2580_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2580_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2579_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx140_2581,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2215_inst_req_0;
      type_cast_2215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2215_inst_req_1;
      type_cast_2215_inst_ack_1<= rack(0);
      type_cast_2215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_2196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2225_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2225_inst_req_0;
      type_cast_2225_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2225_inst_req_1;
      type_cast_2225_inst_ack_1<= rack(0);
      type_cast_2225_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2225_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2193,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_2226,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2235_inst_req_0;
      type_cast_2235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2235_inst_req_1;
      type_cast_2235_inst_ack_1<= rack(0);
      type_cast_2235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2235_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_2199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_2236,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2239_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2239_inst_req_0;
      type_cast_2239_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2239_inst_req_1;
      type_cast_2239_inst_ack_1<= rack(0);
      type_cast_2239_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2239_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_2196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_2240,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2243_inst_req_0;
      type_cast_2243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2243_inst_req_1;
      type_cast_2243_inst_ack_1<= rack(0);
      type_cast_2243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_2208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_2244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2247_inst_req_0;
      type_cast_2247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2247_inst_req_1;
      type_cast_2247_inst_ack_1<= rack(0);
      type_cast_2247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_2205,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_2248,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2256_inst_req_0;
      type_cast_2256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2256_inst_req_1;
      type_cast_2256_inst_ack_1<= rack(0);
      type_cast_2256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_2211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_2257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2260_inst_req_0;
      type_cast_2260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2260_inst_req_1;
      type_cast_2260_inst_ack_1<= rack(0);
      type_cast_2260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_2208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_2261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2270_inst
    process(sext191_2267) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext191_2267(31 downto 0);
      type_cast_2270_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2275_inst
    process(ASHR_i32_i32_2274_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2274_wire(31 downto 0);
      conv90_2276 <= tmp_var; -- 
    end process;
    type_cast_2290_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2290_inst_req_0;
      type_cast_2290_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2290_inst_req_1;
      type_cast_2290_inst_ack_1<= rack(0);
      type_cast_2290_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2290_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2193,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_2291,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2320_inst
    process(sext_2317) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2317(31 downto 0);
      type_cast_2320_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2325_inst
    process(ASHR_i32_i32_2324_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2324_wire(31 downto 0);
      conv108_2326 <= tmp_var; -- 
    end process;
    type_cast_2335_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2335_inst_req_0;
      type_cast_2335_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2335_inst_req_1;
      type_cast_2335_inst_ack_1<= rack(0);
      type_cast_2335_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2335_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_2669,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2335_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2339_inst_req_0;
      type_cast_2339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2339_inst_req_1;
      type_cast_2339_inst_ack_1<= rack(0);
      type_cast_2339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_2676,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2339_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2341_inst_req_0;
      type_cast_2341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2341_inst_req_1;
      type_cast_2341_inst_ack_1<= rack(0);
      type_cast_2341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div11_2232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2341_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2345_inst_req_0;
      type_cast_2345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2345_inst_req_1;
      type_cast_2345_inst_ack_1<= rack(0);
      type_cast_2345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_2682,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2345_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2347_inst_req_0;
      type_cast_2347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2347_inst_req_1;
      type_cast_2347_inst_ack_1<= rack(0);
      type_cast_2347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2347_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2352_inst_req_0;
      type_cast_2352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2352_inst_req_1;
      type_cast_2352_inst_ack_1<= rack(0);
      type_cast_2352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2351_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_2353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2356_inst
    process(conv51_2353) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv51_2353(31 downto 0);
      type_cast_2356_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2358_inst
    process(conv53_2257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv53_2257(31 downto 0);
      type_cast_2358_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2369_inst
    process(conv51_2353) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv51_2353(31 downto 0);
      type_cast_2369_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2371_inst
    process(add_2301) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_2301(31 downto 0);
      type_cast_2371_wire <= tmp_var; -- 
    end process;
    type_cast_2389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2389_inst_req_0;
      type_cast_2389_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2389_inst_req_1;
      type_cast_2389_inst_ack_1<= rack(0);
      type_cast_2389_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2388_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2390,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2393_inst
    process(conv65_2390) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv65_2390(31 downto 0);
      type_cast_2393_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2395_inst
    process(conv53_2257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv53_2257(31 downto 0);
      type_cast_2395_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2406_inst
    process(conv65_2390) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv65_2390(31 downto 0);
      type_cast_2406_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2408_inst
    process(add77_2306) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add77_2306(31 downto 0);
      type_cast_2408_wire <= tmp_var; -- 
    end process;
    type_cast_2426_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2426_inst_req_0;
      type_cast_2426_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2426_inst_req_1;
      type_cast_2426_inst_ack_1<= rack(0);
      type_cast_2426_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2426_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2425_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_2427,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2431_inst_req_0;
      type_cast_2431_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2431_inst_req_1;
      type_cast_2431_inst_ack_1<= rack(0);
      type_cast_2431_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2431_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2430_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_2432,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2455_inst
    process(add94_2452) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add94_2452(31 downto 0);
      type_cast_2455_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2460_inst
    process(ASHR_i32_i32_2459_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2459_wire(31 downto 0);
      shr_2461 <= tmp_var; -- 
    end process;
    type_cast_2465_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2465_inst_req_0;
      type_cast_2465_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2465_inst_req_1;
      type_cast_2465_inst_ack_1<= rack(0);
      type_cast_2465_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2465_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2464_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2466,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2484_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2484_inst_req_0;
      type_cast_2484_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2484_inst_req_1;
      type_cast_2484_inst_ack_1<= rack(0);
      type_cast_2484_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2484_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2483_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_2485,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2538_inst
    process(add115_2515) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add115_2515(31 downto 0);
      type_cast_2538_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2543_inst
    process(ASHR_i32_i32_2542_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2542_wire(31 downto 0);
      shr133_2544 <= tmp_var; -- 
    end process;
    type_cast_2548_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2548_inst_req_0;
      type_cast_2548_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2548_inst_req_1;
      type_cast_2548_inst_ack_1<= rack(0);
      type_cast_2548_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2548_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2547_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom134_2549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2563_inst
    process(add131_2535) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add131_2535(31 downto 0);
      type_cast_2563_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2568_inst
    process(ASHR_i32_i32_2567_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2567_wire(31 downto 0);
      shr138_2569 <= tmp_var; -- 
    end process;
    type_cast_2573_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2573_inst_req_0;
      type_cast_2573_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2573_inst_req_1;
      type_cast_2573_inst_ack_1<= rack(0);
      type_cast_2573_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2573_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2572_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom139_2574,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2591_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2591_inst_req_0;
      type_cast_2591_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2591_inst_req_1;
      type_cast_2591_inst_ack_1<= rack(0);
      type_cast_2591_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2591_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2590_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_2592,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2601_inst
    process(add144_2598) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add144_2598(31 downto 0);
      type_cast_2601_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2603_inst
    process(conv36_2236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv36_2236(31 downto 0);
      type_cast_2603_wire <= tmp_var; -- 
    end process;
    type_cast_2630_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2630_inst_req_0;
      type_cast_2630_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2630_inst_req_1;
      type_cast_2630_inst_ack_1<= rack(0);
      type_cast_2630_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2630_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2629_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv157_2631,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2639_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2639_inst_req_0;
      type_cast_2639_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2639_inst_req_1;
      type_cast_2639_inst_ack_1<= rack(0);
      type_cast_2639_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2639_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp163_2636,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc168_2640,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2655_inst_req_0;
      type_cast_2655_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2655_inst_req_1;
      type_cast_2655_inst_ack_1<= rack(0);
      type_cast_2655_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2654_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_2656,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2672_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2672_inst_req_0;
      type_cast_2672_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2672_inst_req_1;
      type_cast_2672_inst_ack_1<= rack(0);
      type_cast_2672_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2672_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add152_2618,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2672_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2679_inst_req_0;
      type_cast_2679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2679_inst_req_1;
      type_cast_2679_inst_ack_1<= rack(0);
      type_cast_2679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2679_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_2336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2679_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2681_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2681_inst_req_0;
      type_cast_2681_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2681_inst_req_1;
      type_cast_2681_inst_ack_1<= rack(0);
      type_cast_2681_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2681_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc168x_xix_x2_2645,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2681_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2685_inst_req_0;
      type_cast_2685_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2685_inst_req_1;
      type_cast_2685_inst_ack_1<= rack(0);
      type_cast_2685_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2685_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_2342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2685_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2687_inst_req_0;
      type_cast_2687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2687_inst_req_1;
      type_cast_2687_inst_ack_1<= rack(0);
      type_cast_2687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_2651,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2687_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2471_index_1_rename
    process(R_idxprom_2470_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2470_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2470_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2471_index_1_resize
    process(idxprom_2466) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2466;
      ov := iv(13 downto 0);
      R_idxprom_2470_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2471_root_address_inst
    process(array_obj_ref_2471_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2471_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2471_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2554_index_1_rename
    process(R_idxprom134_2553_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom134_2553_resized;
      ov(13 downto 0) := iv;
      R_idxprom134_2553_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2554_index_1_resize
    process(idxprom134_2549) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom134_2549;
      ov := iv(13 downto 0);
      R_idxprom134_2553_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2554_root_address_inst
    process(array_obj_ref_2554_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2554_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2554_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2579_index_1_rename
    process(R_idxprom139_2578_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom139_2578_resized;
      ov(13 downto 0) := iv;
      R_idxprom139_2578_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2579_index_1_resize
    process(idxprom139_2574) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom139_2574;
      ov := iv(13 downto 0);
      R_idxprom139_2578_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2579_root_address_inst
    process(array_obj_ref_2579_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2579_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2579_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2475_addr_0
    process(ptr_deref_2475_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2475_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2475_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2475_base_resize
    process(arrayidx_2473) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2473;
      ov := iv(13 downto 0);
      ptr_deref_2475_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2475_gather_scatter
    process(type_cast_2477_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2477_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2475_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2475_root_address_inst
    process(ptr_deref_2475_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2475_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2475_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2559_addr_0
    process(ptr_deref_2559_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2559_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2559_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2559_base_resize
    process(arrayidx135_2556) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx135_2556;
      ov := iv(13 downto 0);
      ptr_deref_2559_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2559_gather_scatter
    process(ptr_deref_2559_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2559_data_0;
      ov(63 downto 0) := iv;
      tmp136_2560 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2559_root_address_inst
    process(ptr_deref_2559_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2559_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2559_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2583_addr_0
    process(ptr_deref_2583_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2583_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2583_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2583_base_resize
    process(arrayidx140_2581) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx140_2581;
      ov := iv(13 downto 0);
      ptr_deref_2583_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2583_gather_scatter
    process(tmp136_2560) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp136_2560;
      ov(63 downto 0) := iv;
      ptr_deref_2583_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2583_root_address_inst
    process(ptr_deref_2583_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2583_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2583_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2379_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_2378;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2379_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2379_branch_req_0,
          ack0 => if_stmt_2379_branch_ack_0,
          ack1 => if_stmt_2379_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2416_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond192_2415;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2416_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2416_branch_req_0,
          ack0 => if_stmt_2416_branch_ack_0,
          ack1 => if_stmt_2416_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2606_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp147_2605;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2606_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2606_branch_req_0,
          ack0 => if_stmt_2606_branch_ack_0,
          ack1 => if_stmt_2606_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2662_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp178_2661;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2662_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2662_branch_req_0,
          ack0 => if_stmt_2662_branch_ack_0,
          ack1 => if_stmt_2662_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2617_inst
    process(kx_x1_2329) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_2329, type_cast_2616_wire_constant, tmp_var);
      add152_2618 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2625_inst
    process(jx_x1_2342) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_2342, type_cast_2624_wire_constant, tmp_var);
      inc_2626 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2644_inst
    process(inc168_2640, ix_x2_2336) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc168_2640, ix_x2_2336, tmp_var);
      inc168x_xix_x2_2645 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2286_inst
    process(shl_2282, conv38_2240) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_2282, conv38_2240, tmp_var);
      add162_2287 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2295_inst
    process(shl_2282, conv173_2291) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_2282, conv173_2291, tmp_var);
      add177_2296 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2300_inst
    process(conv53_2257, conv173_2291) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv53_2257, conv173_2291, tmp_var);
      add_2301 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2305_inst
    process(conv53_2257, conv38_2240) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv53_2257, conv38_2240, tmp_var);
      add77_2306 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2446_inst
    process(mul93_2442, conv82_2427) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul93_2442, conv82_2427, tmp_var);
      add88_2447 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2451_inst
    process(add88_2447, mul87_2437) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add88_2447, mul87_2437, tmp_var);
      add94_2452 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2509_inst
    process(mul114_2505, conv98_2485) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul114_2505, conv98_2485, tmp_var);
      add106_2510 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2514_inst
    process(add106_2510, mul105_2495) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add106_2510, mul105_2495, tmp_var);
      add115_2515 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2529_inst
    process(mul130_2525, conv98_2485) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul130_2525, conv98_2485, tmp_var);
      add125_2530 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2534_inst
    process(add125_2530, mul124_2520) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add125_2530, mul124_2520, tmp_var);
      add131_2535 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2597_inst
    process(conv143_2592) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv143_2592, type_cast_2596_wire_constant, tmp_var);
      add144_2598 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2377_inst
    process(cmpx_xnot_2366, cmp61_2373) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmpx_xnot_2366, cmp61_2373, tmp_var);
      orx_xcond_2378 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2414_inst
    process(cmp68x_xnot_2403, cmp78_2410) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp68x_xnot_2403, cmp78_2410, tmp_var);
      orx_xcond192_2415 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2274_inst
    process(type_cast_2270_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2270_wire, type_cast_2273_wire_constant, tmp_var);
      ASHR_i32_i32_2274_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2324_inst
    process(type_cast_2320_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2320_wire, type_cast_2323_wire_constant, tmp_var);
      ASHR_i32_i32_2324_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2459_inst
    process(type_cast_2455_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2455_wire, type_cast_2458_wire_constant, tmp_var);
      ASHR_i32_i32_2459_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2542_inst
    process(type_cast_2538_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2538_wire, type_cast_2541_wire_constant, tmp_var);
      ASHR_i32_i32_2542_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2567_inst
    process(type_cast_2563_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2563_wire, type_cast_2566_wire_constant, tmp_var);
      ASHR_i32_i32_2567_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2635_inst
    process(conv157_2631, add162_2287) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv157_2631, add162_2287, tmp_var);
      cmp163_2636 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2660_inst
    process(conv171_2656, add177_2296) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv171_2656, add177_2296, tmp_var);
      cmp178_2661 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2221_inst
    process(conv_2216) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv_2216, type_cast_2220_wire_constant, tmp_var);
      div_2222 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2231_inst
    process(conv10_2226) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv10_2226, type_cast_2230_wire_constant, tmp_var);
      div11_2232 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2252_inst
    process(conv42_2244, conv44_2248) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv42_2244, conv44_2248, tmp_var);
      mul45_2253 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2316_inst
    process(mul_2312, conv36_2236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_2312, conv36_2236, tmp_var);
      sext_2317 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2436_inst
    process(conv86_2432, conv84_2261) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv86_2432, conv84_2261, tmp_var);
      mul87_2437 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2441_inst
    process(conv51_2353, conv90_2276) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv51_2353, conv90_2276, tmp_var);
      mul93_2442 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2494_inst
    process(sub_2490, conv36_2236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_2490, conv36_2236, tmp_var);
      mul105_2495 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2504_inst
    process(sub113_2500, conv108_2326) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub113_2500, conv108_2326, tmp_var);
      mul114_2505 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2519_inst
    process(conv65_2390, conv84_2261) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv65_2390, conv84_2261, tmp_var);
      mul124_2520 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2524_inst
    process(conv51_2353, conv90_2276) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv51_2353, conv90_2276, tmp_var);
      mul130_2525 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2266_inst
    process(mul45_2253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul45_2253, type_cast_2265_wire_constant, tmp_var);
      sext191_2267 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2281_inst
    process(conv53_2257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_2257, type_cast_2280_wire_constant, tmp_var);
      shl_2282 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2311_inst
    process(conv38_2240) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv38_2240, type_cast_2310_wire_constant, tmp_var);
      mul_2312 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2359_inst
    process(type_cast_2356_wire, type_cast_2358_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2356_wire, type_cast_2358_wire, tmp_var);
      cmp_2360 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2372_inst
    process(type_cast_2369_wire, type_cast_2371_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2369_wire, type_cast_2371_wire, tmp_var);
      cmp61_2373 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2396_inst
    process(type_cast_2393_wire, type_cast_2395_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2393_wire, type_cast_2395_wire, tmp_var);
      cmp68_2397 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2409_inst
    process(type_cast_2406_wire, type_cast_2408_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2406_wire, type_cast_2408_wire, tmp_var);
      cmp78_2410 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2604_inst
    process(type_cast_2601_wire, type_cast_2603_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2601_wire, type_cast_2603_wire, tmp_var);
      cmp147_2605 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2489_inst
    process(conv65_2390, conv53_2257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv65_2390, conv53_2257, tmp_var);
      sub_2490 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2499_inst
    process(conv51_2353, conv53_2257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv51_2353, conv53_2257, tmp_var);
      sub113_2500 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_2365_inst
    process(cmp_2360) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp_2360, type_cast_2364_wire_constant, tmp_var);
      cmpx_xnot_2366 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_2402_inst
    process(cmp68_2397) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp68_2397, type_cast_2401_wire_constant, tmp_var);
      cmp68x_xnot_2403 <= tmp_var; --
    end process;
    -- shared split operator group (45) : array_obj_ref_2471_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2470_scaled;
      array_obj_ref_2471_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2471_index_offset_req_0;
      array_obj_ref_2471_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2471_index_offset_req_1;
      array_obj_ref_2471_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : array_obj_ref_2554_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom134_2553_scaled;
      array_obj_ref_2554_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2554_index_offset_req_0;
      array_obj_ref_2554_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2554_index_offset_req_1;
      array_obj_ref_2554_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_2579_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom139_2578_scaled;
      array_obj_ref_2579_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2579_index_offset_req_0;
      array_obj_ref_2579_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2579_index_offset_req_1;
      array_obj_ref_2579_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- unary operator type_cast_2351_inst
    process(ix_x2_2336) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_2336, tmp_var);
      type_cast_2351_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2388_inst
    process(jx_x1_2342) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_2342, tmp_var);
      type_cast_2388_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2425_inst
    process(kx_x1_2329) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2329, tmp_var);
      type_cast_2425_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2430_inst
    process(jx_x1_2342) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_2342, tmp_var);
      type_cast_2430_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2464_inst
    process(shr_2461) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2461, tmp_var);
      type_cast_2464_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2483_inst
    process(kx_x1_2329) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2329, tmp_var);
      type_cast_2483_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2547_inst
    process(shr133_2544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr133_2544, tmp_var);
      type_cast_2547_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2572_inst
    process(shr138_2569) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr138_2569, tmp_var);
      type_cast_2572_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2590_inst
    process(kx_x1_2329) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_2329, tmp_var);
      type_cast_2590_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2629_inst
    process(inc_2626) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2626, tmp_var);
      type_cast_2629_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2654_inst
    process(inc168x_xix_x2_2645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc168x_xix_x2_2645, tmp_var);
      type_cast_2654_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2559_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2559_load_0_req_0;
      ptr_deref_2559_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2559_load_0_req_1;
      ptr_deref_2559_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2559_word_address_0;
      ptr_deref_2559_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2583_store_0 ptr_deref_2475_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2583_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2475_store_0_req_0;
      ptr_deref_2583_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2475_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2583_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2475_store_0_req_1;
      ptr_deref_2583_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2475_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2583_word_address_0 & ptr_deref_2475_word_address_0;
      data_in <= ptr_deref_2583_data_0 & ptr_deref_2475_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_starting_2210_inst RPIPE_Block3_starting_2207_inst RPIPE_Block3_starting_2204_inst RPIPE_Block3_starting_2201_inst RPIPE_Block3_starting_2198_inst RPIPE_Block3_starting_2195_inst RPIPE_Block3_starting_2192_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block3_starting_2210_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_starting_2207_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_starting_2204_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_starting_2201_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_starting_2198_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_starting_2195_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_starting_2192_inst_req_0;
      RPIPE_Block3_starting_2210_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_starting_2207_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_starting_2204_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_starting_2201_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_starting_2198_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_starting_2195_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_starting_2192_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block3_starting_2210_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_starting_2207_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_starting_2204_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_starting_2201_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_starting_2198_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_starting_2195_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_starting_2192_inst_req_1;
      RPIPE_Block3_starting_2210_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_starting_2207_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_starting_2204_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_starting_2201_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_starting_2198_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_starting_2195_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_starting_2192_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call6_2211 <= data_out(55 downto 48);
      call5_2208 <= data_out(47 downto 40);
      call4_2205 <= data_out(39 downto 32);
      call3_2202 <= data_out(31 downto 24);
      call2_2199 <= data_out(23 downto 16);
      call1_2196 <= data_out(15 downto 8);
      call_2193 <= data_out(7 downto 0);
      Block3_starting_read_0_gI: SplitGuardInterface generic map(name => "Block3_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block3_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_starting_pipe_read_req(0),
          oack => Block3_starting_pipe_read_ack(0),
          odata => Block3_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_complete_2692_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_complete_2692_inst_req_0;
      WPIPE_Block3_complete_2692_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_complete_2692_inst_req_1;
      WPIPE_Block3_complete_2692_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2694_wire_constant;
      Block3_complete_write_0_gI: SplitGuardInterface generic map(name => "Block3_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_complete_pipe_write_req(0),
          oack => Block3_complete_pipe_write_ack(0),
          odata => Block3_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(3 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(55 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(255 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(79 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(3 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(7 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_size :  std_logic_vector(31 downto 0);
  signal sendOutput_in_args    : std_logic_vector(31 downto 0);
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_data: std_logic_vector(31 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module zeropad3D
  component zeropad3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block1_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block3_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block1_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block0_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block3_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      Block2_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_data : out  std_logic_vector(31 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D
  signal zeropad3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_start_req : std_logic;
  signal zeropad3D_start_ack : std_logic;
  signal zeropad3D_fin_req   : std_logic;
  signal zeropad3D_fin_ack : std_logic;
  -- declarations related to module zeropad3D_A
  component zeropad3D_A is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block0_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block0_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_A
  signal zeropad3D_A_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_A_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_A_start_req : std_logic;
  signal zeropad3D_A_start_ack : std_logic;
  signal zeropad3D_A_fin_req   : std_logic;
  signal zeropad3D_A_fin_ack : std_logic;
  -- declarations related to module zeropad3D_B
  component zeropad3D_B is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block1_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block1_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_B
  signal zeropad3D_B_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_B_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_B_start_req : std_logic;
  signal zeropad3D_B_start_ack : std_logic;
  signal zeropad3D_B_fin_req   : std_logic;
  signal zeropad3D_B_fin_ack : std_logic;
  -- declarations related to module zeropad3D_C
  component zeropad3D_C is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block2_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_C
  signal zeropad3D_C_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_C_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_C_start_req : std_logic;
  signal zeropad3D_C_start_ack : std_logic;
  signal zeropad3D_C_fin_req   : std_logic;
  signal zeropad3D_C_fin_ack : std_logic;
  -- declarations related to module zeropad3D_D
  component zeropad3D_D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block3_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block3_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_D
  signal zeropad3D_D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_D_start_req : std_logic;
  signal zeropad3D_D_start_ack : std_logic;
  signal zeropad3D_D_fin_req   : std_logic;
  signal zeropad3D_D_fin_ack : std_logic;
  -- aggregate signals for write to pipe Block0_complete
  signal Block0_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block0_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_complete
  signal Block0_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block0_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_starting
  signal Block0_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block0_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_starting
  signal Block0_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block0_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_complete
  signal Block1_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block1_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_complete
  signal Block1_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block1_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_starting
  signal Block1_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block1_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_starting
  signal Block1_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block1_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_complete
  signal Block2_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block2_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_complete
  signal Block2_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block2_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_starting
  signal Block2_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block2_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_starting
  signal Block2_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block2_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_complete
  signal Block3_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block3_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_complete
  signal Block3_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block3_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_starting
  signal Block3_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block3_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_starting
  signal Block3_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block3_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe zeropad_input_pipe
  signal zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe zeropad_output_pipe
  signal zeropad_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal zeropad_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal zeropad_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module sendOutput
  sendOutput_size <= sendOutput_in_args(31 downto 0);
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_data  => sendOutput_call_data,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      call_mdata => sendOutput_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendOutput_size,
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(0 downto 0),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(0 downto 0),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(0 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module zeropad3D
  zeropad3D_instance:zeropad3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_start_req,
      start_ack => zeropad3D_start_ack,
      fin_req => zeropad3D_fin_req,
      fin_ack => zeropad3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      Block0_complete_pipe_read_req => Block0_complete_pipe_read_req(0 downto 0),
      Block0_complete_pipe_read_ack => Block0_complete_pipe_read_ack(0 downto 0),
      Block0_complete_pipe_read_data => Block0_complete_pipe_read_data(7 downto 0),
      Block1_complete_pipe_read_req => Block1_complete_pipe_read_req(0 downto 0),
      Block1_complete_pipe_read_ack => Block1_complete_pipe_read_ack(0 downto 0),
      Block1_complete_pipe_read_data => Block1_complete_pipe_read_data(7 downto 0),
      Block3_complete_pipe_read_req => Block3_complete_pipe_read_req(0 downto 0),
      Block3_complete_pipe_read_ack => Block3_complete_pipe_read_ack(0 downto 0),
      Block3_complete_pipe_read_data => Block3_complete_pipe_read_data(7 downto 0),
      Block2_complete_pipe_read_req => Block2_complete_pipe_read_req(0 downto 0),
      Block2_complete_pipe_read_ack => Block2_complete_pipe_read_ack(0 downto 0),
      Block2_complete_pipe_read_data => Block2_complete_pipe_read_data(7 downto 0),
      zeropad_input_pipe_pipe_read_req => zeropad_input_pipe_pipe_read_req(0 downto 0),
      zeropad_input_pipe_pipe_read_ack => zeropad_input_pipe_pipe_read_ack(0 downto 0),
      zeropad_input_pipe_pipe_read_data => zeropad_input_pipe_pipe_read_data(7 downto 0),
      Block1_starting_pipe_write_req => Block1_starting_pipe_write_req(0 downto 0),
      Block1_starting_pipe_write_ack => Block1_starting_pipe_write_ack(0 downto 0),
      Block1_starting_pipe_write_data => Block1_starting_pipe_write_data(7 downto 0),
      Block0_starting_pipe_write_req => Block0_starting_pipe_write_req(0 downto 0),
      Block0_starting_pipe_write_ack => Block0_starting_pipe_write_ack(0 downto 0),
      Block0_starting_pipe_write_data => Block0_starting_pipe_write_data(7 downto 0),
      Block3_starting_pipe_write_req => Block3_starting_pipe_write_req(0 downto 0),
      Block3_starting_pipe_write_ack => Block3_starting_pipe_write_ack(0 downto 0),
      Block3_starting_pipe_write_data => Block3_starting_pipe_write_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      Block2_starting_pipe_write_req => Block2_starting_pipe_write_req(0 downto 0),
      Block2_starting_pipe_write_ack => Block2_starting_pipe_write_ack(0 downto 0),
      Block2_starting_pipe_write_data => Block2_starting_pipe_write_data(7 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_data => sendOutput_call_data(31 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => zeropad3D_tag_in,
      tag_out => zeropad3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_tag_in <= (others => '0');
  zeropad3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_start_req, start_ack => zeropad3D_start_ack,  fin_req => zeropad3D_fin_req,  fin_ack => zeropad3D_fin_ack);
  -- module zeropad3D_A
  zeropad3D_A_instance:zeropad3D_A-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_A_start_req,
      start_ack => zeropad3D_A_start_ack,
      fin_req => zeropad3D_A_fin_req,
      fin_ack => zeropad3D_A_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_0_sr_req => memory_space_0_sr_req(3 downto 3),
      memory_space_0_sr_ack => memory_space_0_sr_ack(3 downto 3),
      memory_space_0_sr_addr => memory_space_0_sr_addr(55 downto 42),
      memory_space_0_sr_data => memory_space_0_sr_data(255 downto 192),
      memory_space_0_sr_tag => memory_space_0_sr_tag(79 downto 60),
      memory_space_0_sc_req => memory_space_0_sc_req(3 downto 3),
      memory_space_0_sc_ack => memory_space_0_sc_ack(3 downto 3),
      memory_space_0_sc_tag => memory_space_0_sc_tag(7 downto 6),
      Block0_starting_pipe_read_req => Block0_starting_pipe_read_req(0 downto 0),
      Block0_starting_pipe_read_ack => Block0_starting_pipe_read_ack(0 downto 0),
      Block0_starting_pipe_read_data => Block0_starting_pipe_read_data(7 downto 0),
      Block0_complete_pipe_write_req => Block0_complete_pipe_write_req(0 downto 0),
      Block0_complete_pipe_write_ack => Block0_complete_pipe_write_ack(0 downto 0),
      Block0_complete_pipe_write_data => Block0_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_A_tag_in,
      tag_out => zeropad3D_A_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_A_tag_in <= (others => '0');
  zeropad3D_A_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_A_start_req, start_ack => zeropad3D_A_start_ack,  fin_req => zeropad3D_A_fin_req,  fin_ack => zeropad3D_A_fin_ack);
  -- module zeropad3D_B
  zeropad3D_B_instance:zeropad3D_B-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_B_start_req,
      start_ack => zeropad3D_B_start_ack,
      fin_req => zeropad3D_B_fin_req,
      fin_ack => zeropad3D_B_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_0_sr_req => memory_space_0_sr_req(2 downto 2),
      memory_space_0_sr_ack => memory_space_0_sr_ack(2 downto 2),
      memory_space_0_sr_addr => memory_space_0_sr_addr(41 downto 28),
      memory_space_0_sr_data => memory_space_0_sr_data(191 downto 128),
      memory_space_0_sr_tag => memory_space_0_sr_tag(59 downto 40),
      memory_space_0_sc_req => memory_space_0_sc_req(2 downto 2),
      memory_space_0_sc_ack => memory_space_0_sc_ack(2 downto 2),
      memory_space_0_sc_tag => memory_space_0_sc_tag(5 downto 4),
      Block1_starting_pipe_read_req => Block1_starting_pipe_read_req(0 downto 0),
      Block1_starting_pipe_read_ack => Block1_starting_pipe_read_ack(0 downto 0),
      Block1_starting_pipe_read_data => Block1_starting_pipe_read_data(7 downto 0),
      Block1_complete_pipe_write_req => Block1_complete_pipe_write_req(0 downto 0),
      Block1_complete_pipe_write_ack => Block1_complete_pipe_write_ack(0 downto 0),
      Block1_complete_pipe_write_data => Block1_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_B_tag_in,
      tag_out => zeropad3D_B_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_B_tag_in <= (others => '0');
  zeropad3D_B_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_B_start_req, start_ack => zeropad3D_B_start_ack,  fin_req => zeropad3D_B_fin_req,  fin_ack => zeropad3D_B_fin_ack);
  -- module zeropad3D_C
  zeropad3D_C_instance:zeropad3D_C-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_C_start_req,
      start_ack => zeropad3D_C_start_ack,
      fin_req => zeropad3D_C_fin_req,
      fin_ack => zeropad3D_C_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(27 downto 14),
      memory_space_0_sr_data => memory_space_0_sr_data(127 downto 64),
      memory_space_0_sr_tag => memory_space_0_sr_tag(39 downto 20),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 2),
      Block2_starting_pipe_read_req => Block2_starting_pipe_read_req(0 downto 0),
      Block2_starting_pipe_read_ack => Block2_starting_pipe_read_ack(0 downto 0),
      Block2_starting_pipe_read_data => Block2_starting_pipe_read_data(7 downto 0),
      Block2_complete_pipe_write_req => Block2_complete_pipe_write_req(0 downto 0),
      Block2_complete_pipe_write_ack => Block2_complete_pipe_write_ack(0 downto 0),
      Block2_complete_pipe_write_data => Block2_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_C_tag_in,
      tag_out => zeropad3D_C_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_C_tag_in <= (others => '0');
  zeropad3D_C_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_C_start_req, start_ack => zeropad3D_C_start_ack,  fin_req => zeropad3D_C_fin_req,  fin_ack => zeropad3D_C_fin_ack);
  -- module zeropad3D_D
  zeropad3D_D_instance:zeropad3D_D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_D_start_req,
      start_ack => zeropad3D_D_start_ack,
      fin_req => zeropad3D_D_fin_req,
      fin_ack => zeropad3D_D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      Block3_starting_pipe_read_req => Block3_starting_pipe_read_req(0 downto 0),
      Block3_starting_pipe_read_ack => Block3_starting_pipe_read_ack(0 downto 0),
      Block3_starting_pipe_read_data => Block3_starting_pipe_read_data(7 downto 0),
      Block3_complete_pipe_write_req => Block3_complete_pipe_write_req(0 downto 0),
      Block3_complete_pipe_write_ack => Block3_complete_pipe_write_ack(0 downto 0),
      Block3_complete_pipe_write_data => Block3_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_D_tag_in,
      tag_out => zeropad3D_D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_D_tag_in <= (others => '0');
  zeropad3D_D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_D_start_req, start_ack => zeropad3D_D_start_ack,  fin_req => zeropad3D_D_fin_req,  fin_ack => zeropad3D_D_fin_ack);
  Block0_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_complete_pipe_read_req,
      read_ack => Block0_complete_pipe_read_ack,
      read_data => Block0_complete_pipe_read_data,
      write_req => Block0_complete_pipe_write_req,
      write_ack => Block0_complete_pipe_write_ack,
      write_data => Block0_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_starting_pipe_read_req,
      read_ack => Block0_starting_pipe_read_ack,
      read_data => Block0_starting_pipe_read_data,
      write_req => Block0_starting_pipe_write_req,
      write_ack => Block0_starting_pipe_write_ack,
      write_data => Block0_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_complete_pipe_read_req,
      read_ack => Block1_complete_pipe_read_ack,
      read_data => Block1_complete_pipe_read_data,
      write_req => Block1_complete_pipe_write_req,
      write_ack => Block1_complete_pipe_write_ack,
      write_data => Block1_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_starting_pipe_read_req,
      read_ack => Block1_starting_pipe_read_ack,
      read_data => Block1_starting_pipe_read_data,
      write_req => Block1_starting_pipe_write_req,
      write_ack => Block1_starting_pipe_write_ack,
      write_data => Block1_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_complete_pipe_read_req,
      read_ack => Block2_complete_pipe_read_ack,
      read_data => Block2_complete_pipe_read_data,
      write_req => Block2_complete_pipe_write_req,
      write_ack => Block2_complete_pipe_write_ack,
      write_data => Block2_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_starting_pipe_read_req,
      read_ack => Block2_starting_pipe_read_ack,
      read_data => Block2_starting_pipe_read_data,
      write_req => Block2_starting_pipe_write_req,
      write_ack => Block2_starting_pipe_write_ack,
      write_data => Block2_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_complete_pipe_read_req,
      read_ack => Block3_complete_pipe_read_ack,
      read_data => Block3_complete_pipe_read_data,
      write_req => Block3_complete_pipe_write_req,
      write_ack => Block3_complete_pipe_write_ack,
      write_data => Block3_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_starting_pipe_read_req,
      read_ack => Block3_starting_pipe_read_ack,
      read_data => Block3_starting_pipe_read_data,
      write_req => Block3_starting_pipe_write_req,
      write_ack => Block3_starting_pipe_write_ack,
      write_data => Block3_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_input_pipe_pipe_read_req,
      read_ack => zeropad_input_pipe_pipe_read_ack,
      read_data => zeropad_input_pipe_pipe_read_data,
      write_req => zeropad_input_pipe_pipe_write_req,
      write_ack => zeropad_input_pipe_pipe_write_ack,
      write_data => zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_output_pipe_pipe_read_req,
      read_ack => zeropad_output_pipe_pipe_read_ack,
      read_data => zeropad_output_pipe_pipe_read_data,
      write_req => zeropad_output_pipe_pipe_write_req,
      write_ack => zeropad_output_pipe_pipe_write_ack,
      write_data => zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 4,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyROM_memory_space_2: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
