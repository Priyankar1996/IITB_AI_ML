-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package baud_control_calculator_global_package is -- 
  component baud_control_calculator is -- 
    port (-- 
      clk : in std_logic;
      reset : in std_logic); -- 
    -- 
  end component;
  -- 
end package baud_control_calculator_global_package;
