-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity fill_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(63 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity fill_T;
architecture fill_T_arch of fill_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(63 downto 0);
  signal addr_update_enable: Boolean;
  -- output port buffer signals
  signal fill_T_CP_0_start: Boolean;
  signal fill_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_41_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_41_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_41_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_41_inst_ack_1 : boolean;
  signal CONCAT_u240_u256_48_inst_req_0 : boolean;
  signal CONCAT_u240_u256_48_inst_ack_0 : boolean;
  signal CONCAT_u240_u256_48_inst_req_1 : boolean;
  signal CONCAT_u240_u256_48_inst_ack_1 : boolean;
  signal addr_of_63_final_reg_req_0 : boolean;
  signal addr_of_63_final_reg_ack_0 : boolean;
  signal addr_of_63_final_reg_req_1 : boolean;
  signal addr_of_63_final_reg_ack_1 : boolean;
  signal if_stmt_50_branch_req_0 : boolean;
  signal if_stmt_50_branch_ack_1 : boolean;
  signal if_stmt_50_branch_ack_0 : boolean;
  signal phi_stmt_23_req_0 : boolean;
  signal phi_stmt_29_req_0 : boolean;
  signal nmycount_39_28_buf_req_0 : boolean;
  signal nmycount_39_28_buf_ack_0 : boolean;
  signal nmycount_39_28_buf_req_1 : boolean;
  signal nmycount_39_28_buf_ack_1 : boolean;
  signal phi_stmt_23_req_1 : boolean;
  signal ninput_word_49_33_buf_req_0 : boolean;
  signal ninput_word_49_33_buf_ack_0 : boolean;
  signal ninput_word_49_33_buf_req_1 : boolean;
  signal ninput_word_49_33_buf_ack_1 : boolean;
  signal phi_stmt_29_req_1 : boolean;
  signal phi_stmt_23_ack_0 : boolean;
  signal phi_stmt_29_ack_0 : boolean;
  signal array_obj_ref_62_index_offset_req_0 : boolean;
  signal array_obj_ref_62_index_offset_ack_0 : boolean;
  signal array_obj_ref_62_index_offset_req_1 : boolean;
  signal array_obj_ref_62_index_offset_ack_1 : boolean;
  signal ptr_deref_66_store_0_req_0 : boolean;
  signal ptr_deref_66_store_0_ack_0 : boolean;
  signal ptr_deref_66_store_0_req_1 : boolean;
  signal ptr_deref_66_store_0_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "fill_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  fill_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "fill_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= fill_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,fill_T_CP_0_start,"fill_T cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,fill_T_CP_0_symbol, "fill_T cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  fill_T_CP_0: Block -- control-path 
    signal fill_T_CP_0_elements: BooleanArray(29 downto 0);
    -- 
  begin -- 
    fill_T_CP_0_elements(0) <= fill_T_CP_0_start;
    fill_T_CP_0_symbol <= fill_T_CP_0_elements(29);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	8 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_21/$entry
      -- CP-element group 0: 	 branch_block_stmt_21/branch_block_stmt_21__entry__
      -- CP-element group 0: 	 branch_block_stmt_21/merge_stmt_22__entry__
      -- CP-element group 0: 	 branch_block_stmt_21/merge_stmt_22_dead_link/$entry
      -- 
    -- logger for CP element group fill_T_CP_0_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	22 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	5 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_21/merge_stmt_22__exit__
      -- CP-element group 1: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49__entry__
      -- CP-element group 1: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/$entry
      -- CP-element group 1: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_update_start_
      -- CP-element group 1: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_Update/cr
      -- 
    -- logger for CP element group fill_T_CP_0_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:RPIPE_maxpool_input_pipe_41_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:CONCAT_u240_u256_48_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_24_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_24_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => RPIPE_maxpool_input_pipe_41_inst_req_0); -- 
    cr_43_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_43_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => CONCAT_u240_u256_48_inst_req_1); -- 
    fill_T_CP_0_elements(1) <= fill_T_CP_0_elements(22);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_update_start_
      -- CP-element group 2: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_Update/cr
      -- 
    -- logger for CP element group fill_T_CP_0_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:RPIPE_maxpool_input_pipe_41_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:RPIPE_maxpool_input_pipe_41_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_25_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_41_inst_ack_0, ack => fill_T_CP_0_elements(2)); -- 
    cr_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(2), ack => RPIPE_maxpool_input_pipe_41_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/RPIPE_maxpool_input_pipe_41_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_Sample/rr
      -- 
    -- logger for CP element group fill_T_CP_0_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:RPIPE_maxpool_input_pipe_41_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:CONCAT_u240_u256_48_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_30_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_41_inst_ack_1, ack => fill_T_CP_0_elements(3)); -- 
    rr_38_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_38_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(3), ack => CONCAT_u240_u256_48_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_Sample/ra
      -- 
    -- logger for CP element group fill_T_CP_0_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:CONCAT_u240_u256_48_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_39_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u240_u256_48_inst_ack_0, ack => fill_T_CP_0_elements(4)); -- 
    -- CP-element group 5:  branch  transition  place  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (27) 
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/$entry
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/$exit
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/ULT_u4_u1_53_inputs/$entry
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/ULT_u4_u1_53_inputs/$exit
      -- CP-element group 5: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49__exit__
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50__entry__
      -- CP-element group 5: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/$exit
      -- CP-element group 5: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_21/assign_stmt_39_to_assign_stmt_49/CONCAT_u240_u256_48_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_dead_link/$entry
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/$entry
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/$exit
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/SplitProtocol/$exit
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/SplitProtocol/Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/SplitProtocol/Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/SplitProtocol/Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/ULT_u4_u1_53/SplitProtocol/Update/ca
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_eval_test/branch_req
      -- CP-element group 5: 	 branch_block_stmt_21/ULT_u4_u1_53_place
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_if_link/$entry
      -- CP-element group 5: 	 branch_block_stmt_21/if_stmt_50_else_link/$entry
      -- 
    -- logger for CP element group fill_T_CP_0_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:CONCAT_u240_u256_48_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:if_stmt_50_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_44_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u240_u256_48_inst_ack_1, ack => fill_T_CP_0_elements(5)); -- 
    branch_req_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(5), ack => if_stmt_50_branch_req_0); -- 
    -- CP-element group 6:  fork  transition  place  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	16 
    -- CP-element group 6: 	15 
    -- CP-element group 6: 	12 
    -- CP-element group 6: 	13 
    -- CP-element group 6:  members (18) 
      -- CP-element group 6: 	 branch_block_stmt_21/if_stmt_50_if_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_21/if_stmt_50_if_link/if_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_21/loopback
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/req
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/req
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/Interlock/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/Interlock/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/Interlock/Sample/req
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/Interlock/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/Interlock/Update/req
      -- 
    -- logger for CP element group fill_T_CP_0_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:if_stmt_50_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:nmycount_39_28_buf_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:nmycount_39_28_buf_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:ninput_word_49_33_buf_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:ninput_word_49_33_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_76_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_50_branch_ack_1, ack => fill_T_CP_0_elements(6)); -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(6), ack => nmycount_39_28_buf_req_0); -- 
    req_125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(6), ack => nmycount_39_28_buf_req_1); -- 
    req_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(6), ack => ninput_word_49_33_buf_req_0); -- 
    req_145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(6), ack => ninput_word_49_33_buf_req_1); -- 
    -- CP-element group 7:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	23 
    -- CP-element group 7: 	24 
    -- CP-element group 7: 	26 
    -- CP-element group 7: 	28 
    -- CP-element group 7:  members (30) 
      -- CP-element group 7: 	 branch_block_stmt_21/$exit
      -- CP-element group 7: 	 branch_block_stmt_21/branch_block_stmt_21__exit__
      -- CP-element group 7: 	 branch_block_stmt_21/if_stmt_50__exit__
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/$entry
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/req
      -- CP-element group 7: 	 branch_block_stmt_21/if_stmt_50_else_link/$exit
      -- CP-element group 7: 	 branch_block_stmt_21/if_stmt_50_else_link/else_choice_transition
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/$entry
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_update_start_
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resized_1
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scaled_1
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_computed_1
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/$entry
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/$exit
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/index_resize_req
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/index_resize_ack
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/$entry
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/$exit
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/scale_rename_req
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/scale_rename_ack
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_update_start
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/$entry
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/req
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/$entry
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/req
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_update_start_
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/$entry
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/$entry
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/$entry
      -- CP-element group 7: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group fill_T_CP_0_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:if_stmt_50_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:addr_of_63_final_reg_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:array_obj_ref_62_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:array_obj_ref_62_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:ptr_deref_66_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_80_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_50_branch_ack_0, ack => fill_T_CP_0_elements(7)); -- 
    req_201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(7), ack => addr_of_63_final_reg_req_1); -- 
    req_181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(7), ack => array_obj_ref_62_index_offset_req_0); -- 
    req_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(7), ack => array_obj_ref_62_index_offset_req_1); -- 
    cr_251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(7), ack => ptr_deref_66_store_0_req_1); -- 
    -- CP-element group 8:  fork  transition  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_23/$entry
      -- CP-element group 8: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_29/$entry
      -- CP-element group 8: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_29/phi_stmt_29_sources/$entry
      -- 
    -- logger for CP element group fill_T_CP_0_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    fill_T_CP_0_elements(8) <= fill_T_CP_0_elements(0);
    -- CP-element group 9:  transition  output  delay-element  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_23/$exit
      -- CP-element group 9: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/$exit
      -- CP-element group 9: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/type_cast_27_konst_delay_trans
      -- CP-element group 9: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_23/phi_stmt_23_req
      -- 
    -- logger for CP element group fill_T_CP_0_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:phi_stmt_23_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_23_req_96_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_23_req_96_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(9), ack => phi_stmt_23_req_0); -- 
    -- Element group fill_T_CP_0_elements(9) is a control-delay.
    cp_element_9_delay: control_delay_element  generic map(name => " 9_delay", delay_value => 1)  port map(req => fill_T_CP_0_elements(8), ack => fill_T_CP_0_elements(9), clk => clk, reset =>reset);
    -- CP-element group 10:  transition  output  delay-element  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (4) 
      -- CP-element group 10: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_29/$exit
      -- CP-element group 10: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_29/phi_stmt_29_sources/$exit
      -- CP-element group 10: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_29/phi_stmt_29_sources/type_cast_32_konst_delay_trans
      -- CP-element group 10: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/phi_stmt_29/phi_stmt_29_req
      -- 
    -- logger for CP element group fill_T_CP_0_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:phi_stmt_29_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_29_req_104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_29_req_104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => phi_stmt_29_req_0); -- 
    -- Element group fill_T_CP_0_elements(10) is a control-delay.
    cp_element_10_delay: control_delay_element  generic map(name => " 10_delay", delay_value => 1)  port map(req => fill_T_CP_0_elements(8), ack => fill_T_CP_0_elements(10), clk => clk, reset =>reset);
    -- CP-element group 11:  join  transition  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	19 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_21/merge_stmt_22__entry___PhiReq/$exit
      -- 
    -- logger for CP element group fill_T_CP_0_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    fill_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(9) & fill_T_CP_0_elements(10);
      gj_fill_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	6 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/ack
      -- 
    -- logger for CP element group fill_T_CP_0_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:nmycount_39_28_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_39_28_buf_ack_0, ack => fill_T_CP_0_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	6 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/ack
      -- 
    -- logger for CP element group fill_T_CP_0_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:nmycount_39_28_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_39_28_buf_ack_1, ack => fill_T_CP_0_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	18 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/$exit
      -- CP-element group 14: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/$exit
      -- CP-element group 14: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/$exit
      -- CP-element group 14: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_23/phi_stmt_23_req
      -- 
    -- logger for CP element group fill_T_CP_0_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:phi_stmt_23_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_23_req_127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_23_req_127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(14), ack => phi_stmt_23_req_1); -- 
    fill_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(12) & fill_T_CP_0_elements(13);
      gj_fill_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	6 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/Interlock/Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/Interlock/Sample/ack
      -- 
    -- logger for CP element group fill_T_CP_0_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:ninput_word_49_33_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_49_33_buf_ack_0, ack => fill_T_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	6 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/Interlock/Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/Interlock/Update/ack
      -- 
    -- logger for CP element group fill_T_CP_0_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:ninput_word_49_33_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_49_33_buf_ack_1, ack => fill_T_CP_0_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/$exit
      -- CP-element group 17: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/$exit
      -- CP-element group 17: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_sources/Interlock/$exit
      -- CP-element group 17: 	 branch_block_stmt_21/loopback_PhiReq/phi_stmt_29/phi_stmt_29_req
      -- 
    -- logger for CP element group fill_T_CP_0_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:phi_stmt_29_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_29_req_147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_29_req_147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(17), ack => phi_stmt_29_req_1); -- 
    fill_T_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(16) & fill_T_CP_0_elements(15);
      gj_fill_T_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: 	14 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_21/loopback_PhiReq/$exit
      -- 
    -- logger for CP element group fill_T_CP_0_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    fill_T_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(17) & fill_T_CP_0_elements(14);
      gj_fill_T_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  merge  fork  transition  place  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: 	11 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_21/merge_stmt_22_PhiReqMerge
      -- CP-element group 19: 	 branch_block_stmt_21/merge_stmt_22_PhiAck/$entry
      -- 
    -- logger for CP element group fill_T_CP_0_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    fill_T_CP_0_elements(19) <= OrReduce(fill_T_CP_0_elements(18) & fill_T_CP_0_elements(11));
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_21/merge_stmt_22_PhiAck/phi_stmt_23_ack
      -- 
    -- logger for CP element group fill_T_CP_0_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:phi_stmt_23_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_23_ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_23_ack_0, ack => fill_T_CP_0_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_21/merge_stmt_22_PhiAck/phi_stmt_29_ack
      -- 
    -- logger for CP element group fill_T_CP_0_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:phi_stmt_29_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_29_ack_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_29_ack_0, ack => fill_T_CP_0_elements(21)); -- 
    -- CP-element group 22:  join  transition  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	1 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_21/merge_stmt_22_PhiAck/$exit
      -- 
    -- logger for CP element group fill_T_CP_0_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    fill_T_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(20) & fill_T_CP_0_elements(21);
      gj_fill_T_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	7 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	29 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_sample_complete
      -- CP-element group 23: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/$exit
      -- CP-element group 23: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group fill_T_CP_0_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:array_obj_ref_62_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_index_offset_ack_0, ack => fill_T_CP_0_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	7 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (11) 
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/$entry
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/req
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_sample_start_
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_root_address_calculated
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_offset_calculated
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/$exit
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/ack
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/$entry
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/$exit
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/sum_rename_req
      -- CP-element group 24: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/sum_rename_ack
      -- 
    -- logger for CP element group fill_T_CP_0_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:array_obj_ref_62_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:addr_of_63_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_index_offset_ack_1, ack => fill_T_CP_0_elements(24)); -- 
    req_196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(24), ack => addr_of_63_final_reg_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/$exit
      -- CP-element group 25: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/ack
      -- CP-element group 25: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_sample_completed_
      -- 
    -- logger for CP element group fill_T_CP_0_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:addr_of_63_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_63_final_reg_ack_0, ack => fill_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	7 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (28) 
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/$exit
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/ack
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_update_completed_
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_sample_start_
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_address_calculated
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_address_calculated
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_root_address_calculated
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_address_resized
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/$entry
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/$exit
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/base_resize_req
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/base_resize_ack
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/$entry
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/$exit
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/sum_rename_req
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/sum_rename_ack
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/$entry
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/$exit
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/root_register_req
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/root_register_ack
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/$entry
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/$entry
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/$exit
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/split_req
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/split_ack
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/$entry
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/$entry
      -- CP-element group 26: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group fill_T_CP_0_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:addr_of_63_final_reg_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:ptr_deref_66_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_63_final_reg_ack_1, ack => fill_T_CP_0_elements(26)); -- 
    rr_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(26), ack => ptr_deref_66_store_0_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_sample_completed_
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/$exit
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/$exit
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group fill_T_CP_0_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:ptr_deref_66_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_66_store_0_ack_0, ack => fill_T_CP_0_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	7 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (5) 
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_update_completed_
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/$exit
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/$exit
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group fill_T_CP_0_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:ptr_deref_66_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_66_store_0_ack_1, ack => fill_T_CP_0_elements(28)); -- 
    -- CP-element group 29:  join  transition  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 $exit
      -- CP-element group 29: 	 assign_stmt_64_to_assign_stmt_68/$exit
      -- 
    -- logger for CP element group fill_T_CP_0_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and fill_T_CP_0_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:fill_T:CP:fill_T_CP_0_elements(29) fired."); 
        -- 
      end if; --
    end process; 
    fill_T_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(23) & fill_T_CP_0_elements(28);
      gj_fill_T_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(29), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_addr_61_resized : std_logic_vector(13 downto 0);
    signal R_addr_61_scaled : std_logic_vector(13 downto 0);
    signal ULT_u4_u1_53_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_62_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_62_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_62_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_62_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_62_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_62_root_address : std_logic_vector(13 downto 0);
    signal input_word_29 : std_logic_vector(255 downto 0);
    signal konst_37_wire_constant : std_logic_vector(3 downto 0);
    signal konst_52_wire_constant : std_logic_vector(3 downto 0);
    signal mycount_23 : std_logic_vector(3 downto 0);
    signal ninput_word_49 : std_logic_vector(255 downto 0);
    signal ninput_word_49_33_buffered : std_logic_vector(255 downto 0);
    signal nmycount_39 : std_logic_vector(3 downto 0);
    signal nmycount_39_28_buffered : std_logic_vector(3 downto 0);
    signal ptr_64 : std_logic_vector(31 downto 0);
    signal ptr_deref_66_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_66_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_66_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_66_wire : std_logic_vector(255 downto 0);
    signal ptr_deref_66_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_66_word_offset_0 : std_logic_vector(13 downto 0);
    signal slice_46_wire : std_logic_vector(239 downto 0);
    signal type_cast_27_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_32_wire_constant : std_logic_vector(255 downto 0);
    signal val_42 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_62_constant_part_of_offset <= "00000000000000";
    array_obj_ref_62_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_62_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_62_resized_base_address <= "00000000000000";
    konst_37_wire_constant <= "0001";
    konst_52_wire_constant <= "1111";
    ptr_deref_66_word_offset_0 <= "00000000000000";
    type_cast_27_wire_constant <= "0000";
    type_cast_32_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    -- logger for phi phi_stmt_23
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_23_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:fill_T:DP:phi_stmt_23:input-0 type_cast_27_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_27_wire_constant));
          --
        end if;
        if phi_stmt_23_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:fill_T:DP:phi_stmt_23:input-1 nmycount_39_28_buffered= " & Convert_SLV_To_Hex_String(nmycount_39_28_buffered));
          --
        end if;
        if phi_stmt_23_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:fill_T:DP:phi_stmt_23:sample-completed");
          --
        end if;
        if phi_stmt_23_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:fill_T:DP:phi_stmt_23:output mycount_23= " & Convert_SLV_To_Hex_String(mycount_23));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_23: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_27_wire_constant & nmycount_39_28_buffered;
      req <= phi_stmt_23_req_0 & phi_stmt_23_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_23",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_23_ack_0,
          idata => idata,
          odata => mycount_23,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_23
    -- logger for phi phi_stmt_29
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_29_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:fill_T:DP:phi_stmt_29:input-0 type_cast_32_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_32_wire_constant));
          --
        end if;
        if phi_stmt_29_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:fill_T:DP:phi_stmt_29:input-1 ninput_word_49_33_buffered= " & Convert_SLV_To_Hex_String(ninput_word_49_33_buffered));
          --
        end if;
        if phi_stmt_29_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:fill_T:DP:phi_stmt_29:sample-completed");
          --
        end if;
        if phi_stmt_29_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:fill_T:DP:phi_stmt_29:output input_word_29= " & Convert_SLV_To_Hex_String(input_word_29));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_29: Block -- phi operator 
      signal idata: std_logic_vector(511 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_32_wire_constant & ninput_word_49_33_buffered;
      req <= phi_stmt_29_req_0 & phi_stmt_29_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_29",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 256) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_29_ack_0,
          idata => idata,
          odata => input_word_29,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_29
    -- logger for split-operator slice_46_inst flow-through 
    process(slice_46_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:slice_46_inst:flowthrough inputs: " & " input_word_29 = "& Convert_SLV_To_Hex_String(input_word_29) & " outputs:" & " slice_46_wire= "  & Convert_SLV_To_Hex_String(slice_46_wire));
      --
    end process; 
    -- flow-through slice operator slice_46_inst
    slice_46_wire <= input_word_29(239 downto 0);
    -- logger for split-operator addr_of_63_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_63_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:addr_of_63_final_reg:started:   inputs: " & " array_obj_ref_62_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_62_root_address));
          --
        end if; 
        if addr_of_63_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:addr_of_63_final_reg:finished:  outputs: " & " ptr_64= "  & Convert_SLV_To_Hex_String(ptr_64));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_63_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_63_final_reg_req_0;
      addr_of_63_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_63_final_reg_req_1;
      addr_of_63_final_reg_ack_1<= rack(0);
      addr_of_63_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_63_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_62_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator ninput_word_49_33_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ninput_word_49_33_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:ninput_word_49_33_buf:started:   inputs: " & " ninput_word_49 = "& Convert_SLV_To_Hex_String(ninput_word_49));
          --
        end if; 
        if ninput_word_49_33_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:ninput_word_49_33_buf:finished:  outputs: " & " ninput_word_49_33_buffered= "  & Convert_SLV_To_Hex_String(ninput_word_49_33_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    ninput_word_49_33_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ninput_word_49_33_buf_req_0;
      ninput_word_49_33_buf_ack_0<= wack(0);
      rreq(0) <= ninput_word_49_33_buf_req_1;
      ninput_word_49_33_buf_ack_1<= rack(0);
      ninput_word_49_33_buf : InterlockBuffer generic map ( -- 
        name => "ninput_word_49_33_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 256,
        out_data_width => 256,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ninput_word_49,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ninput_word_49_33_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator nmycount_39_28_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if nmycount_39_28_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:nmycount_39_28_buf:started:   inputs: " & " nmycount_39 = "& Convert_SLV_To_Hex_String(nmycount_39));
          --
        end if; 
        if nmycount_39_28_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:nmycount_39_28_buf:finished:  outputs: " & " nmycount_39_28_buffered= "  & Convert_SLV_To_Hex_String(nmycount_39_28_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    nmycount_39_28_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_39_28_buf_req_0;
      nmycount_39_28_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_39_28_buf_req_1;
      nmycount_39_28_buf_ack_1<= rack(0);
      nmycount_39_28_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_39_28_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_39,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_39_28_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_62_index_1_rename flow-through 
    process(R_addr_61_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:array_obj_ref_62_index_1_rename:flowthrough  inputs: " & " R_addr_61_resized = "& Convert_SLV_To_Hex_String(R_addr_61_resized) & "outputs: " & " R_addr_61_scaled= "  & Convert_SLV_To_Hex_String(R_addr_61_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_62_index_1_rename
    process(R_addr_61_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_61_resized;
      ov(13 downto 0) := iv;
      R_addr_61_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_62_index_1_resize flow-through 
    process(R_addr_61_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:array_obj_ref_62_index_1_resize:flowthrough  inputs: " & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & "outputs: " & " R_addr_61_resized= "  & Convert_SLV_To_Hex_String(R_addr_61_resized));
      --
    end process; 
    -- equivalence array_obj_ref_62_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(13 downto 0);
      R_addr_61_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_62_root_address_inst flow-through 
    process(array_obj_ref_62_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:array_obj_ref_62_root_address_inst:flowthrough  inputs: " & " array_obj_ref_62_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_62_final_offset) & "outputs: " & " array_obj_ref_62_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_62_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_62_root_address_inst
    process(array_obj_ref_62_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_62_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_62_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_66_addr_0 flow-through 
    process(ptr_deref_66_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:ptr_deref_66_addr_0:flowthrough  inputs: " & " ptr_deref_66_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_66_root_address) & "outputs: " & " ptr_deref_66_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_66_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_66_addr_0
    process(ptr_deref_66_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_66_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_66_base_resize flow-through 
    process(ptr_deref_66_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:ptr_deref_66_base_resize:flowthrough  inputs: " & " ptr_64 = "& Convert_SLV_To_Hex_String(ptr_64) & "outputs: " & " ptr_deref_66_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_66_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_66_base_resize
    process(ptr_64) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_64;
      ov := iv(13 downto 0);
      ptr_deref_66_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_66_gather_scatter flow-through 
    process(ptr_deref_66_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:ptr_deref_66_gather_scatter:flowthrough  inputs: " & " ninput_word_49 = "& Convert_SLV_To_Hex_String(ninput_word_49) & "outputs: " & " ptr_deref_66_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_66_data_0));
      --
    end process; 
    -- equivalence ptr_deref_66_gather_scatter
    process(ninput_word_49) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ninput_word_49;
      ov(255 downto 0) := iv;
      ptr_deref_66_data_0 <= ov(255 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_66_root_address_inst flow-through 
    process(ptr_deref_66_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:ptr_deref_66_root_address_inst:flowthrough  inputs: " & " ptr_deref_66_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_66_resized_base_address) & "outputs: " & " ptr_deref_66_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_66_root_address));
      --
    end process; 
    -- equivalence ptr_deref_66_root_address_inst
    process(ptr_deref_66_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_66_root_address <= ov(13 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_50_branch_req_0," req0 if_stmt_50_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_50_branch_ack_0," ack0 if_stmt_50_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_50_branch_ack_1," ack1 if_stmt_50_branch");
    if_stmt_50_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u4_u1_53_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_50_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_50_branch_req_0,
          ack0 => if_stmt_50_branch_ack_0,
          ack1 => if_stmt_50_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u4_u4_38_inst flow-through 
    process(nmycount_39) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:ADD_u4_u4_38_inst:flowthrough inputs: " & " mycount_23 = "& Convert_SLV_To_Hex_String(mycount_23) & " konst_37_wire_constant = "& Convert_SLV_To_Hex_String(konst_37_wire_constant) & " outputs:" & " nmycount_39= "  & Convert_SLV_To_Hex_String(nmycount_39));
      --
    end process; 
    -- binary operator ADD_u4_u4_38_inst
    process(mycount_23) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_23, konst_37_wire_constant, tmp_var);
      nmycount_39 <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u240_u256_48_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u240_u256_48_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:CONCAT_u240_u256_48_inst:started:   inputs: " & " slice_46_wire = "& Convert_SLV_To_Hex_String(slice_46_wire) & " val_42 = "& Convert_SLV_To_Hex_String(val_42));
          --
        end if; 
        if CONCAT_u240_u256_48_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:CONCAT_u240_u256_48_inst:finished:  outputs: " & " ninput_word_49= "  & Convert_SLV_To_Hex_String(ninput_word_49));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (1) : CONCAT_u240_u256_48_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(255 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_46_wire & val_42;
      ninput_word_49 <= data_out(255 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u240_u256_48_inst_req_0;
      CONCAT_u240_u256_48_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u240_u256_48_inst_req_1;
      CONCAT_u240_u256_48_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 240,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 256,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- logger for split-operator ULT_u4_u1_53_inst flow-through 
    process(ULT_u4_u1_53_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:ULT_u4_u1_53_inst:flowthrough inputs: " & " mycount_23 = "& Convert_SLV_To_Hex_String(mycount_23) & " konst_52_wire_constant = "& Convert_SLV_To_Hex_String(konst_52_wire_constant) & " outputs:" & " ULT_u4_u1_53_wire= "  & Convert_SLV_To_Hex_String(ULT_u4_u1_53_wire));
      --
    end process; 
    -- binary operator ULT_u4_u1_53_inst
    process(mycount_23) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_23, konst_52_wire_constant, tmp_var);
      ULT_u4_u1_53_wire <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_62_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_62_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:array_obj_ref_62_index_offset:started:   inputs: " & " R_addr_61_scaled = "& Convert_SLV_To_Hex_String(R_addr_61_scaled) & " array_obj_ref_62_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_62_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_62_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:array_obj_ref_62_index_offset:finished:  outputs: " & " array_obj_ref_62_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_62_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (3) : array_obj_ref_62_index_offset 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_61_scaled;
      array_obj_ref_62_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_62_index_offset_req_0;
      array_obj_ref_62_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_62_index_offset_req_1;
      array_obj_ref_62_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- logger for split-operator ptr_deref_66_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_66_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:ptr_deref_66_store_0:started:   inputs: " & " ptr_deref_66_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_66_word_address_0) & " ptr_deref_66_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_66_data_0));
          --
        end if; 
        if ptr_deref_66_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:ptr_deref_66_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_66_store_0_req_0,
      ptr_deref_66_store_0_ack_0,
      ptr_deref_66_store_0_req_1,
      ptr_deref_66_store_0_ack_1,
      "ptr_deref_66_store_0",
      "memory_space_1" ,
      ptr_deref_66_data_0,
      ptr_deref_66_word_address_0,
      "ptr_deref_66_data_0",
      "ptr_deref_66_word_address_0" -- 
    );
    -- shared store operator group (0) : ptr_deref_66_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_66_store_0_req_0;
      ptr_deref_66_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_66_store_0_req_1;
      ptr_deref_66_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_66_word_address_0;
      data_in <= ptr_deref_66_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 256,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(255 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logger for split-operator RPIPE_maxpool_input_pipe_41_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_41_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:RPIPE_maxpool_input_pipe_41_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_41_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:fill_T:DP:RPIPE_maxpool_input_pipe_41_inst:finished:  outputs: " & " val_42= "  & Convert_SLV_To_Hex_String(val_42));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_41_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_41_inst_req_0;
      RPIPE_maxpool_input_pipe_41_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_41_inst_req_1;
      RPIPE_maxpool_input_pipe_41_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      val_42 <= data_out(15 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end fill_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(8 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_call_acks : in   std_logic_vector(0 downto 0);
    maxPool4_call_data : out  std_logic_vector(159 downto 0);
    maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
    maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_return_acks : in   std_logic_vector(0 downto 0);
    maxPool4_return_data : in   std_logic_vector(7 downto 0);
    maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
    sendB_call_reqs : out  std_logic_vector(0 downto 0);
    sendB_call_acks : in   std_logic_vector(0 downto 0);
    sendB_call_tag  :  out  std_logic_vector(0 downto 0);
    sendB_return_reqs : out  std_logic_vector(0 downto 0);
    sendB_return_acks : in   std_logic_vector(0 downto 0);
    sendB_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool3D;
architecture maxPool3D_arch of maxPool3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal maxPool3D_CP_4436_start: Boolean;
  signal maxPool3D_CP_4436_symbol: Boolean;
  -- volatile/operator module components. 
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(8 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      fill_T_call_reqs : out  std_logic_vector(0 downto 0);
      fill_T_call_acks : in   std_logic_vector(0 downto 0);
      fill_T_call_data : out  std_logic_vector(63 downto 0);
      fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
      fill_T_return_reqs : out  std_logic_vector(0 downto 0);
      fill_T_return_acks : in   std_logic_vector(0 downto 0);
      fill_T_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      output : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1712_call_req_0 : boolean;
  signal W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_ack_0 : boolean;
  signal type_cast_1852_inst_req_1 : boolean;
  signal type_cast_1852_inst_ack_1 : boolean;
  signal type_cast_1948_inst_req_1 : boolean;
  signal if_stmt_2023_branch_req_0 : boolean;
  signal W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_req_0 : boolean;
  signal type_cast_1852_inst_ack_0 : boolean;
  signal call_stmt_1939_call_req_0 : boolean;
  signal call_stmt_1712_call_ack_1 : boolean;
  signal call_stmt_1712_call_ack_0 : boolean;
  signal call_stmt_1712_call_req_1 : boolean;
  signal W_rowx_x1_1974_delayed_4_0_1990_inst_req_0 : boolean;
  signal type_cast_1979_inst_ack_0 : boolean;
  signal do_while_stmt_1842_branch_ack_0 : boolean;
  signal type_cast_1957_inst_ack_1 : boolean;
  signal type_cast_2031_inst_ack_1 : boolean;
  signal type_cast_1979_inst_req_0 : boolean;
  signal type_cast_2031_inst_req_1 : boolean;
  signal W_rowx_x1_1974_delayed_4_0_1990_inst_ack_1 : boolean;
  signal call_stmt_1939_call_ack_0 : boolean;
  signal type_cast_1948_inst_ack_1 : boolean;
  signal call_stmt_1939_call_req_1 : boolean;
  signal type_cast_2031_inst_ack_0 : boolean;
  signal type_cast_1957_inst_req_1 : boolean;
  signal W_rowx_x1_1974_delayed_4_0_1990_inst_req_1 : boolean;
  signal type_cast_2031_inst_req_0 : boolean;
  signal type_cast_1979_inst_ack_1 : boolean;
  signal type_cast_1979_inst_req_1 : boolean;
  signal type_cast_1988_inst_req_0 : boolean;
  signal type_cast_1988_inst_ack_0 : boolean;
  signal type_cast_2010_inst_ack_1 : boolean;
  signal do_while_stmt_1842_branch_ack_1 : boolean;
  signal W_rowx_x1_1974_delayed_4_0_1990_inst_ack_0 : boolean;
  signal type_cast_1988_inst_req_1 : boolean;
  signal W_colx_x1_1949_delayed_2_0_1959_inst_req_0 : boolean;
  signal W_colx_x1_1949_delayed_2_0_1959_inst_ack_0 : boolean;
  signal type_cast_1957_inst_req_0 : boolean;
  signal type_cast_2010_inst_req_1 : boolean;
  signal type_cast_1862_inst_req_0 : boolean;
  signal type_cast_1988_inst_ack_1 : boolean;
  signal type_cast_1948_inst_req_0 : boolean;
  signal type_cast_1957_inst_ack_0 : boolean;
  signal phi_stmt_1854_req_1 : boolean;
  signal type_cast_1948_inst_ack_0 : boolean;
  signal if_stmt_2023_branch_ack_1 : boolean;
  signal W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_req_1 : boolean;
  signal W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_ack_1 : boolean;
  signal call_stmt_1939_call_ack_1 : boolean;
  signal type_cast_1852_inst_req_0 : boolean;
  signal type_cast_1858_inst_ack_1 : boolean;
  signal type_cast_1858_inst_req_1 : boolean;
  signal ptr_deref_1724_load_0_req_0 : boolean;
  signal ptr_deref_1724_load_0_ack_0 : boolean;
  signal ptr_deref_1724_load_0_req_1 : boolean;
  signal ptr_deref_1724_load_0_ack_1 : boolean;
  signal type_cast_1870_inst_ack_1 : boolean;
  signal W_inc_1956_delayed_1_0_1967_inst_ack_1 : boolean;
  signal type_cast_1870_inst_req_1 : boolean;
  signal type_cast_1870_inst_ack_0 : boolean;
  signal type_cast_1870_inst_req_0 : boolean;
  signal W_inc_1956_delayed_1_0_1967_inst_req_1 : boolean;
  signal type_cast_1858_inst_ack_0 : boolean;
  signal ptr_deref_1736_load_0_req_0 : boolean;
  signal type_cast_1866_inst_ack_1 : boolean;
  signal ptr_deref_1736_load_0_ack_0 : boolean;
  signal type_cast_1858_inst_req_0 : boolean;
  signal ptr_deref_1736_load_0_req_1 : boolean;
  signal type_cast_1866_inst_req_1 : boolean;
  signal ptr_deref_1736_load_0_ack_1 : boolean;
  signal W_inc_1956_delayed_1_0_1967_inst_ack_0 : boolean;
  signal type_cast_2010_inst_ack_0 : boolean;
  signal type_cast_1866_inst_ack_0 : boolean;
  signal type_cast_1866_inst_req_0 : boolean;
  signal W_inc_1956_delayed_1_0_1967_inst_req_0 : boolean;
  signal phi_stmt_1854_ack_0 : boolean;
  signal phi_stmt_1854_req_0 : boolean;
  signal ptr_deref_1748_addr_0_req_0 : boolean;
  signal ptr_deref_1748_addr_0_ack_0 : boolean;
  signal ptr_deref_1748_addr_0_req_1 : boolean;
  signal ptr_deref_1748_addr_0_ack_1 : boolean;
  signal ptr_deref_1748_addr_1_req_0 : boolean;
  signal ptr_deref_1748_addr_1_ack_0 : boolean;
  signal ptr_deref_1748_addr_1_req_1 : boolean;
  signal ptr_deref_1748_addr_1_ack_1 : boolean;
  signal type_cast_2010_inst_req_0 : boolean;
  signal if_stmt_2023_branch_ack_0 : boolean;
  signal ptr_deref_1748_addr_2_req_0 : boolean;
  signal ptr_deref_1748_addr_2_ack_0 : boolean;
  signal ptr_deref_1748_addr_2_req_1 : boolean;
  signal W_colx_x1_1949_delayed_2_0_1959_inst_ack_1 : boolean;
  signal ptr_deref_1748_addr_2_ack_1 : boolean;
  signal type_cast_1862_inst_ack_1 : boolean;
  signal type_cast_1862_inst_req_1 : boolean;
  signal ptr_deref_1748_addr_3_req_0 : boolean;
  signal W_colx_x1_1949_delayed_2_0_1959_inst_req_1 : boolean;
  signal ptr_deref_1748_addr_3_ack_0 : boolean;
  signal ptr_deref_1748_addr_3_req_1 : boolean;
  signal ptr_deref_1748_addr_3_ack_1 : boolean;
  signal ptr_deref_1748_load_0_req_0 : boolean;
  signal ptr_deref_1748_load_0_ack_0 : boolean;
  signal type_cast_1862_inst_ack_0 : boolean;
  signal ptr_deref_1748_load_1_req_0 : boolean;
  signal ptr_deref_1748_load_1_ack_0 : boolean;
  signal ptr_deref_1748_load_2_req_0 : boolean;
  signal ptr_deref_1748_load_2_ack_0 : boolean;
  signal ptr_deref_1748_load_3_req_0 : boolean;
  signal ptr_deref_1748_load_3_ack_0 : boolean;
  signal ptr_deref_1748_load_0_req_1 : boolean;
  signal ptr_deref_1748_load_0_ack_1 : boolean;
  signal ptr_deref_1748_load_1_req_1 : boolean;
  signal ptr_deref_1748_load_1_ack_1 : boolean;
  signal ptr_deref_1748_load_2_req_1 : boolean;
  signal ptr_deref_1748_load_2_ack_1 : boolean;
  signal ptr_deref_1748_load_3_req_1 : boolean;
  signal ptr_deref_1748_load_3_ack_1 : boolean;
  signal ptr_deref_1760_load_0_req_0 : boolean;
  signal ptr_deref_1760_load_0_ack_0 : boolean;
  signal ptr_deref_1760_load_0_req_1 : boolean;
  signal ptr_deref_1760_load_0_ack_1 : boolean;
  signal call_stmt_1787_call_req_0 : boolean;
  signal call_stmt_1787_call_ack_0 : boolean;
  signal call_stmt_1787_call_req_1 : boolean;
  signal call_stmt_1787_call_ack_1 : boolean;
  signal do_while_stmt_1842_branch_req_0 : boolean;
  signal phi_stmt_1844_req_0 : boolean;
  signal phi_stmt_1844_req_1 : boolean;
  signal phi_stmt_1844_ack_0 : boolean;
  signal type_cast_1847_inst_req_0 : boolean;
  signal type_cast_1847_inst_ack_0 : boolean;
  signal type_cast_1847_inst_req_1 : boolean;
  signal type_cast_1847_inst_ack_1 : boolean;
  signal phi_stmt_1849_req_0 : boolean;
  signal phi_stmt_1849_req_1 : boolean;
  signal phi_stmt_1849_ack_0 : boolean;
  signal call_stmt_2035_call_req_0 : boolean;
  signal call_stmt_2035_call_ack_0 : boolean;
  signal call_stmt_2035_call_req_1 : boolean;
  signal call_stmt_2035_call_ack_1 : boolean;
  signal type_cast_2039_inst_req_0 : boolean;
  signal type_cast_2039_inst_ack_0 : boolean;
  signal type_cast_2039_inst_req_1 : boolean;
  signal type_cast_2039_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_2046_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_2046_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_2046_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_2046_inst_ack_1 : boolean;
  signal call_stmt_2050_call_req_0 : boolean;
  signal call_stmt_2050_call_ack_0 : boolean;
  signal call_stmt_2050_call_req_1 : boolean;
  signal call_stmt_2050_call_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool3D_CP_4436_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool3D_CP_4436_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool3D_CP_4436_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool3D_CP_4436_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,maxPool3D_CP_4436_start,"maxPool3D cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,maxPool3D_CP_4436_symbol, "maxPool3D cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool3D_CP_4436: Block -- control-path 
    signal maxPool3D_CP_4436_elements: BooleanArray(176 downto 0);
    -- 
  begin -- 
    maxPool3D_CP_4436_elements(0) <= maxPool3D_CP_4436_start;
    maxPool3D_CP_4436_symbol <= maxPool3D_CP_4436_elements(176);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_1711/call_stmt_1712__entry__
      -- CP-element group 0: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1711/$entry
      -- CP-element group 0: 	 branch_block_stmt_1711/call_stmt_1712/$entry
      -- CP-element group 0: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_Update/ccr
      -- CP-element group 0: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1711/branch_block_stmt_1711__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1712_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1712_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_4478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(0), ack => call_stmt_1712_call_req_0); -- 
    ccr_4483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(0), ack => call_stmt_1712_call_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	164 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	165 
    -- CP-element group 1: 	166 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_1711/do_while_stmt_1842__exit__
      -- CP-element group 1: 	 branch_block_stmt_1711/if_stmt_2023_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_1711/R_whilex_xbody_whilex_xend_taken_2024_place
      -- CP-element group 1: 	 branch_block_stmt_1711/if_stmt_2023_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1711/if_stmt_2023_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_1711/if_stmt_2023_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1711/if_stmt_2023__entry__
      -- CP-element group 1: 	 branch_block_stmt_1711/if_stmt_2023_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_1711/if_stmt_2023_else_link/$entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:if_stmt_2023_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_5128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(1), ack => if_stmt_2023_branch_req_0); -- 
    maxPool3D_CP_4436_elements(1) <= maxPool3D_CP_4436_elements(164);
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_Sample/cra
      -- CP-element group 2: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_sample_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1712_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_4479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1712_call_ack_0, ack => maxPool3D_CP_4436_elements(2)); -- 
    -- CP-element group 3:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	5 
    -- CP-element group 3: 	6 
    -- CP-element group 3: 	7 
    -- CP-element group 3: 	8 
    -- CP-element group 3: 	11 
    -- CP-element group 3: 	12 
    -- CP-element group 3: 	13 
    -- CP-element group 3: 	14 
    -- CP-element group 3: 	15 
    -- CP-element group 3: 	16 
    -- CP-element group 3: 	17 
    -- CP-element group 3: 	18 
    -- CP-element group 3: 	24 
    -- CP-element group 3: 	25 
    -- CP-element group 3: 	26 
    -- CP-element group 3: 	27 
    -- CP-element group 3: 	29 
    -- CP-element group 3: 	30 
    -- CP-element group 3:  members (125) 
      -- CP-element group 3: 	 branch_block_stmt_1711/call_stmt_1712__exit__
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_Update/cca
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1711/call_stmt_1712/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_1711/call_stmt_1712/call_stmt_1712_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784__entry__
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_sample_start
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_update_start
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_0_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_0_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_0_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_0_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_1_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_1_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_1_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_1_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_2_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_2_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_2_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_2_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_3_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_3_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_3_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_3_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_0/cr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_1/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_1/cr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_2/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_2/cr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_3/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_3/cr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_base_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_word_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_root_address_calculated
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_base_address_resized
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_base_addr_resize/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_base_addr_resize/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_base_addr_resize/base_resize_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_base_addr_resize/base_resize_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_base_plus_offset/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_base_plus_offset/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_base_plus_offset/sum_rename_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_base_plus_offset/sum_rename_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_word_addrgen/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_word_addrgen/$exit
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_word_addrgen/root_register_req
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_word_addrgen/root_register_ack
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/word_access_complete/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/word_access_complete/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1712_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1724_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1724_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1736_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1736_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_3_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1760_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1760_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_4484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1712_call_ack_1, ack => maxPool3D_CP_4436_elements(3)); -- 
    rr_4520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1724_load_0_req_0); -- 
    cr_4531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1724_load_0_req_1); -- 
    rr_4570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1736_load_0_req_0); -- 
    cr_4581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1736_load_0_req_1); -- 
    rr_4613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_addr_0_req_0); -- 
    cr_4618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_addr_0_req_1); -- 
    rr_4623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_addr_1_req_0); -- 
    cr_4628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_addr_1_req_1); -- 
    rr_4633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_addr_2_req_0); -- 
    cr_4638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_addr_2_req_1); -- 
    rr_4643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_addr_3_req_0); -- 
    cr_4648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_addr_3_req_1); -- 
    cr_4685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_load_0_req_1); -- 
    cr_4690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_load_1_req_1); -- 
    cr_4695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_load_2_req_1); -- 
    cr_4700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1748_load_3_req_1); -- 
    rr_4739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1760_load_0_req_0); -- 
    cr_4750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(3), ack => ptr_deref_1760_load_0_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Sample/word_access_start/$exit
      -- CP-element group 4: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1724_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1724_load_0_ack_0, ack => maxPool3D_CP_4436_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	3 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	31 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/word_access_complete/$exit
      -- CP-element group 5: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/word_access_complete/word_0/ca
      -- CP-element group 5: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/ptr_deref_1724_Merge/$entry
      -- CP-element group 5: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/ptr_deref_1724_Merge/$exit
      -- CP-element group 5: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/ptr_deref_1724_Merge/merge_req
      -- CP-element group 5: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1724_Update/ptr_deref_1724_Merge/merge_ack
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1724_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1724_load_0_ack_1, ack => maxPool3D_CP_4436_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1736_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1736_load_0_ack_0, ack => maxPool3D_CP_4436_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	3 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	31 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/word_access_complete/word_0/ca
      -- CP-element group 7: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/ptr_deref_1736_Merge/$entry
      -- CP-element group 7: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/ptr_deref_1736_Merge/$exit
      -- CP-element group 7: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/ptr_deref_1736_Merge/merge_req
      -- CP-element group 7: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1736_Update/ptr_deref_1736_Merge/merge_ack
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1736_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1736_load_0_ack_1, ack => maxPool3D_CP_4436_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	3 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	19 
    -- CP-element group 8: 	20 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	22 
    -- CP-element group 8:  members (11) 
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_0/rr
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_1/$entry
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_1/rr
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_2/$entry
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_2/rr
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_3/$entry
      -- CP-element group 8: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_3/rr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_3_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(8), ack => ptr_deref_1748_load_0_req_0); -- 
    rr_4664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(8), ack => ptr_deref_1748_load_1_req_0); -- 
    rr_4669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(8), ack => ptr_deref_1748_load_2_req_0); -- 
    rr_4674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(8), ack => ptr_deref_1748_load_3_req_0); -- 
    maxPool3D_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool3D_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(3) & maxPool3D_CP_4436_elements(10);
      gj_maxPool3D_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	17 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	31 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_sample_complete
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "maxPool3D_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(11) & maxPool3D_CP_4436_elements(13) & maxPool3D_CP_4436_elements(15) & maxPool3D_CP_4436_elements(17);
      gj_maxPool3D_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	18 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_update_complete
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(10) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(12) & maxPool3D_CP_4436_elements(14) & maxPool3D_CP_4436_elements(16) & maxPool3D_CP_4436_elements(18);
      gj_maxPool3D_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	3 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_0_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_0_Sample/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_addr_0_ack_0, ack => maxPool3D_CP_4436_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	3 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_0_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_0_Update/ca
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_addr_0_ack_1, ack => maxPool3D_CP_4436_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	9 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_1_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_1_Sample/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_addr_1_ack_0, ack => maxPool3D_CP_4436_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	3 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_1_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_1_Update/ca
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_addr_1_ack_1, ack => maxPool3D_CP_4436_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	3 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	9 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_2_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_2_Sample/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_addr_2_ack_0, ack => maxPool3D_CP_4436_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	3 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	10 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_2_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_2_Update/ca
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_addr_2_ack_1, ack => maxPool3D_CP_4436_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	9 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_3_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_3_Sample/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_addr_3_ack_0, ack => maxPool3D_CP_4436_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	3 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	10 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_3_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_word_addrgen_3_Update/ca
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_addr_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_addr_3_ack_1, ack => maxPool3D_CP_4436_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	8 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	23 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_load_0_ack_0, ack => maxPool3D_CP_4436_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	8 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	23 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_1/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_load_1_ack_0, ack => maxPool3D_CP_4436_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_2/$exit
      -- CP-element group 21: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_2/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_load_2_ack_0, ack => maxPool3D_CP_4436_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	8 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_3/$exit
      -- CP-element group 22: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/word_3/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_load_3_ack_0, ack => maxPool3D_CP_4436_elements(22)); -- 
    -- CP-element group 23:  join  transition  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: 	20 
    -- CP-element group 23: 	21 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(19) & maxPool3D_CP_4436_elements(20) & maxPool3D_CP_4436_elements(21) & maxPool3D_CP_4436_elements(22);
      gj_maxPool3D_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	3 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	28 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_load_0_ack_1, ack => maxPool3D_CP_4436_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	3 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_1/$exit
      -- CP-element group 25: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_1/ca
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_load_1_ack_1, ack => maxPool3D_CP_4436_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	3 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_2/$exit
      -- CP-element group 26: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_2/ca
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_load_2_ack_1, ack => maxPool3D_CP_4436_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	3 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_3/$exit
      -- CP-element group 27: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/word_3/ca
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1748_load_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1748_load_3_ack_1, ack => maxPool3D_CP_4436_elements(27)); -- 
    -- CP-element group 28:  join  transition  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: 	25 
    -- CP-element group 28: 	26 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (7) 
      -- CP-element group 28: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/ptr_deref_1748_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/ptr_deref_1748_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/ptr_deref_1748_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1748_Update/ptr_deref_1748_Merge/merge_ack
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(24) & maxPool3D_CP_4436_elements(25) & maxPool3D_CP_4436_elements(26) & maxPool3D_CP_4436_elements(27);
      gj_maxPool3D_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	3 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1760_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1760_load_0_ack_0, ack => maxPool3D_CP_4436_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	3 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/ptr_deref_1760_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/ptr_deref_1760_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/ptr_deref_1760_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/ptr_deref_1760_Update/ptr_deref_1760_Merge/merge_ack
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:ptr_deref_1760_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1760_load_0_ack_1, ack => maxPool3D_CP_4436_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	5 
    -- CP-element group 31: 	7 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (10) 
      -- CP-element group 31: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784/$exit
      -- CP-element group 31: 	 branch_block_stmt_1711/call_stmt_1787__entry__
      -- CP-element group 31: 	 branch_block_stmt_1711/assign_stmt_1721_to_assign_stmt_1784__exit__
      -- CP-element group 31: 	 branch_block_stmt_1711/call_stmt_1787/$entry
      -- CP-element group 31: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_Sample/crr
      -- CP-element group 31: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_Update/ccr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1787_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1787_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_4767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(31), ack => call_stmt_1787_call_req_0); -- 
    ccr_4772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(31), ack => call_stmt_1787_call_req_1); -- 
    maxPool3D_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(5) & maxPool3D_CP_4436_elements(7) & maxPool3D_CP_4436_elements(9) & maxPool3D_CP_4436_elements(28) & maxPool3D_CP_4436_elements(30);
      gj_maxPool3D_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_Sample/cra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1787_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_4768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1787_call_ack_0, ack => maxPool3D_CP_4436_elements(32)); -- 
    -- CP-element group 33:  transition  place  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (17) 
      -- CP-element group 33: 	 branch_block_stmt_1711/do_while_stmt_1842__entry__
      -- CP-element group 33: 	 branch_block_stmt_1711/entry_whilex_xbody
      -- CP-element group 33: 	 branch_block_stmt_1711/assign_stmt_1794_to_assign_stmt_1823__entry__
      -- CP-element group 33: 	 branch_block_stmt_1711/call_stmt_1787__exit__
      -- CP-element group 33: 	 branch_block_stmt_1711/merge_stmt_1825__exit__
      -- CP-element group 33: 	 branch_block_stmt_1711/assign_stmt_1794_to_assign_stmt_1823__exit__
      -- CP-element group 33: 	 branch_block_stmt_1711/call_stmt_1787/$exit
      -- CP-element group 33: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1711/call_stmt_1787/call_stmt_1787_Update/cca
      -- CP-element group 33: 	 branch_block_stmt_1711/assign_stmt_1794_to_assign_stmt_1823/$entry
      -- CP-element group 33: 	 branch_block_stmt_1711/assign_stmt_1794_to_assign_stmt_1823/$exit
      -- CP-element group 33: 	 branch_block_stmt_1711/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_1711/entry_whilex_xbody_PhiReq/$exit
      -- CP-element group 33: 	 branch_block_stmt_1711/merge_stmt_1825_PhiReqMerge
      -- CP-element group 33: 	 branch_block_stmt_1711/merge_stmt_1825_PhiAck/$entry
      -- CP-element group 33: 	 branch_block_stmt_1711/merge_stmt_1825_PhiAck/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1787_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_4773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1787_call_ack_1, ack => maxPool3D_CP_4436_elements(33)); -- 
    -- CP-element group 34:  transition  place  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_1711/do_while_stmt_1842/$entry
      -- CP-element group 34: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842__entry__
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(34) <= maxPool3D_CP_4436_elements(33);
    -- CP-element group 35:  merge  place  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	164 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842__exit__
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(35) is bound as output of CP function.
    -- CP-element group 36:  merge  place  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	39 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1711/do_while_stmt_1842/loop_back
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(36) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(36) is bound as output of CP function.
    -- CP-element group 37:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	42 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	162 
    -- CP-element group 37: 	163 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1711/do_while_stmt_1842/loop_taken/$entry
      -- CP-element group 37: 	 branch_block_stmt_1711/do_while_stmt_1842/loop_exit/$entry
      -- CP-element group 37: 	 branch_block_stmt_1711/do_while_stmt_1842/condition_done
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(37) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(37) <= maxPool3D_CP_4436_elements(42);
    -- CP-element group 38:  branch  place  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	161 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1711/do_while_stmt_1842/loop_body_done
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(38) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(38) <= maxPool3D_CP_4436_elements(161);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	36 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	51 
    -- CP-element group 39: 	72 
    -- CP-element group 39: 	93 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(39) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(39) <= maxPool3D_CP_4436_elements(36);
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	53 
    -- CP-element group 40: 	74 
    -- CP-element group 40: 	95 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(40) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(40) <= maxPool3D_CP_4436_elements(34);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	47 
    -- CP-element group 41: 	48 
    -- CP-element group 41: 	66 
    -- CP-element group 41: 	67 
    -- CP-element group 41: 	87 
    -- CP-element group 41: 	88 
    -- CP-element group 41: 	160 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/$entry
      -- CP-element group 41: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/loop_body_start
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(41) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	46 
    -- CP-element group 42: 	159 
    -- CP-element group 42: 	160 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	37 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/condition_evaluated
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:do_while_stmt_1842_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_4791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(42), ack => do_while_stmt_1842_branch_req_0); -- 
    maxPool3D_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(46) & maxPool3D_CP_4436_elements(159) & maxPool3D_CP_4436_elements(160);
      gj_maxPool3D_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	47 
    -- CP-element group 43: 	66 
    -- CP-element group 43: 	87 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	46 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	68 
    -- CP-element group 43: 	89 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/aggregated_phi_sample_req
      -- CP-element group 43: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_sample_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(43) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(47) & maxPool3D_CP_4436_elements(66) & maxPool3D_CP_4436_elements(87) & maxPool3D_CP_4436_elements(46);
      gj_maxPool3D_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	49 
    -- CP-element group 44: 	69 
    -- CP-element group 44: 	90 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	125 
    -- CP-element group 44: 	137 
    -- CP-element group 44: 	141 
    -- CP-element group 44: 	145 
    -- CP-element group 44: 	149 
    -- CP-element group 44: 	153 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44: 	66 
    -- CP-element group 44: 	87 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/aggregated_phi_sample_ack
      -- CP-element group 44: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_sample_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(44) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(49) & maxPool3D_CP_4436_elements(69) & maxPool3D_CP_4436_elements(90);
      gj_maxPool3D_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	48 
    -- CP-element group 45: 	67 
    -- CP-element group 45: 	88 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	70 
    -- CP-element group 45: 	91 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/aggregated_phi_update_req
      -- CP-element group 45: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_update_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(45) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(48) & maxPool3D_CP_4436_elements(67) & maxPool3D_CP_4436_elements(88);
      gj_maxPool3D_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	50 
    -- CP-element group 46: 	71 
    -- CP-element group 46: 	92 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	42 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	43 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(50) & maxPool3D_CP_4436_elements(71) & maxPool3D_CP_4436_elements(92);
      gj_maxPool3D_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	41 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	147 
    -- CP-element group 47: 	151 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	43 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(47) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(41) & maxPool3D_CP_4436_elements(44) & maxPool3D_CP_4436_elements(147) & maxPool3D_CP_4436_elements(151);
      gj_maxPool3D_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	41 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: 	118 
    -- CP-element group 48: 	150 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	45 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(48) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(41) & maxPool3D_CP_4436_elements(50) & maxPool3D_CP_4436_elements(118) & maxPool3D_CP_4436_elements(150);
      gj_maxPool3D_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	44 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_sample_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(49) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(49) is bound as output of CP function.
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	46 
    -- CP-element group 50: 	116 
    -- CP-element group 50: 	148 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_update_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(50) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(50) is bound as output of CP function.
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	39 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_loopback_trigger
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(51) <= maxPool3D_CP_4436_elements(39);
    -- CP-element group 52:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (2) 
      -- CP-element group 52: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_loopback_sample_req
      -- CP-element group 52: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_loopback_sample_req_ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:phi_stmt_1844_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1844_loopback_sample_req_4806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1844_loopback_sample_req_4806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(52), ack => phi_stmt_1844_req_0); -- 
    -- Element group maxPool3D_CP_4436_elements(52) is bound as output of CP function.
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	40 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_entry_trigger
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(53) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(53) <= maxPool3D_CP_4436_elements(40);
    -- CP-element group 54:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_entry_sample_req
      -- CP-element group 54: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_entry_sample_req_ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:phi_stmt_1844_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1844_entry_sample_req_4809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1844_entry_sample_req_4809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(54), ack => phi_stmt_1844_req_1); -- 
    -- Element group maxPool3D_CP_4436_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_phi_mux_ack
      -- CP-element group 55: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1844_phi_mux_ack_ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:phi_stmt_1844_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1844_phi_mux_ack_4812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1844_ack_0, ack => maxPool3D_CP_4436_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_sample_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(56) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_update_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(57) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_Sample/rr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1847_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(58), ack => type_cast_1847_inst_req_0); -- 
    maxPool3D_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(56) & maxPool3D_CP_4436_elements(60);
      gj_maxPool3D_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_update_start_
      -- CP-element group 59: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_Update/cr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1847_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(59), ack => type_cast_1847_inst_req_1); -- 
    maxPool3D_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(57) & maxPool3D_CP_4436_elements(61);
      gj_maxPool3D_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (4) 
      -- CP-element group 60: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_sample_completed__ps
      -- CP-element group 60: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_Sample/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1847_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1847_inst_ack_0, ack => maxPool3D_CP_4436_elements(60)); -- 
    -- CP-element group 61:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_update_completed__ps
      -- CP-element group 61: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1847_Update/ca
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1847_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1847_inst_ack_1, ack => maxPool3D_CP_4436_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_rowx_x1_at_entry_1848_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_rowx_x1_at_entry_1848_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_rowx_x1_at_entry_1848_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_rowx_x1_at_entry_1848_sample_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(62) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_rowx_x1_at_entry_1848_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_rowx_x1_at_entry_1848_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(63) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_rowx_x1_at_entry_1848_update_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(64) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(64) <= maxPool3D_CP_4436_elements(65);
    -- CP-element group 65:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	64 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_rowx_x1_at_entry_1848_update_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(65) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => maxPool3D_CP_4436_elements(63), ack => maxPool3D_CP_4436_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  join  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	41 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	44 
    -- CP-element group 66: 	143 
    -- CP-element group 66: 	155 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	43 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(66) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(41) & maxPool3D_CP_4436_elements(44) & maxPool3D_CP_4436_elements(143) & maxPool3D_CP_4436_elements(155);
      gj_maxPool3D_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	41 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	71 
    -- CP-element group 67: 	114 
    -- CP-element group 67: 	134 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	45 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(67) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(41) & maxPool3D_CP_4436_elements(71) & maxPool3D_CP_4436_elements(114) & maxPool3D_CP_4436_elements(134);
      gj_maxPool3D_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	43 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_sample_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(68) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(68) <= maxPool3D_CP_4436_elements(43);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	44 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_sample_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(69) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(69) is bound as output of CP function.
    -- CP-element group 70:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	45 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_update_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(70) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(70) <= maxPool3D_CP_4436_elements(45);
    -- CP-element group 71:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	46 
    -- CP-element group 71: 	112 
    -- CP-element group 71: 	132 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	67 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_update_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(71) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(71) is bound as output of CP function.
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	39 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_loopback_trigger
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(72) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(72) <= maxPool3D_CP_4436_elements(39);
    -- CP-element group 73:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_loopback_sample_req
      -- CP-element group 73: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_loopback_sample_req_ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:phi_stmt_1849_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1849_loopback_sample_req_4850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1849_loopback_sample_req_4850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(73), ack => phi_stmt_1849_req_0); -- 
    -- Element group maxPool3D_CP_4436_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	40 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_entry_trigger
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(74) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(74) <= maxPool3D_CP_4436_elements(40);
    -- CP-element group 75:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_entry_sample_req
      -- CP-element group 75: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_entry_sample_req_ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:phi_stmt_1849_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1849_entry_sample_req_4853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1849_entry_sample_req_4853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(75), ack => phi_stmt_1849_req_1); -- 
    -- Element group maxPool3D_CP_4436_elements(75) is bound as output of CP function.
    -- CP-element group 76:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_phi_mux_ack
      -- CP-element group 76: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1849_phi_mux_ack_ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:phi_stmt_1849_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1849_phi_mux_ack_4856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1849_ack_0, ack => maxPool3D_CP_4436_elements(76)); -- 
    -- CP-element group 77:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_sample_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(77) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_update_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(78) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(78) is bound as output of CP function.
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	81 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1852_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(79), ack => type_cast_1852_inst_req_0); -- 
    maxPool3D_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(77) & maxPool3D_CP_4436_elements(81);
      gj_maxPool3D_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1852_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(80), ack => type_cast_1852_inst_req_1); -- 
    maxPool3D_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(78) & maxPool3D_CP_4436_elements(82);
      gj_maxPool3D_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	79 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_sample_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1852_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1852_inst_ack_0, ack => maxPool3D_CP_4436_elements(81)); -- 
    -- CP-element group 82:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1852_update_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1852_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1852_inst_ack_1, ack => maxPool3D_CP_4436_elements(82)); -- 
    -- CP-element group 83:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_colx_x1_at_entry_1853_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_colx_x1_at_entry_1853_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_colx_x1_at_entry_1853_sample_completed__ps
      -- CP-element group 83: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_colx_x1_at_entry_1853_sample_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(83) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_colx_x1_at_entry_1853_update_start_
      -- CP-element group 84: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_colx_x1_at_entry_1853_update_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(84) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(84) is bound as output of CP function.
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_colx_x1_at_entry_1853_update_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(85) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(85) <= maxPool3D_CP_4436_elements(86);
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	85 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_colx_x1_at_entry_1853_update_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(86) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => maxPool3D_CP_4436_elements(84), ack => maxPool3D_CP_4436_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	41 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	44 
    -- CP-element group 87: 	127 
    -- CP-element group 87: 	139 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	43 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(87) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(41) & maxPool3D_CP_4436_elements(44) & maxPool3D_CP_4436_elements(127) & maxPool3D_CP_4436_elements(139);
      gj_maxPool3D_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	41 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	92 
    -- CP-element group 88: 	110 
    -- CP-element group 88: 	126 
    -- CP-element group 88: 	138 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	45 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(88) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(41) & maxPool3D_CP_4436_elements(92) & maxPool3D_CP_4436_elements(110) & maxPool3D_CP_4436_elements(126) & maxPool3D_CP_4436_elements(138);
      gj_maxPool3D_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	43 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_sample_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(89) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(89) <= maxPool3D_CP_4436_elements(43);
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	44 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_sample_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(90) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(90) is bound as output of CP function.
    -- CP-element group 91:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	45 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_update_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(91) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(91) <= maxPool3D_CP_4436_elements(45);
    -- CP-element group 92:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	46 
    -- CP-element group 92: 	108 
    -- CP-element group 92: 	124 
    -- CP-element group 92: 	136 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	88 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_update_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_update_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(92) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(92) is bound as output of CP function.
    -- CP-element group 93:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	39 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_loopback_trigger
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(93) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(93) <= maxPool3D_CP_4436_elements(39);
    -- CP-element group 94:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_loopback_sample_req
      -- CP-element group 94: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_loopback_sample_req_ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:phi_stmt_1854_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1854_loopback_sample_req_4894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1854_loopback_sample_req_4894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(94), ack => phi_stmt_1854_req_1); -- 
    -- Element group maxPool3D_CP_4436_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	40 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_entry_trigger
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(95) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(95) <= maxPool3D_CP_4436_elements(40);
    -- CP-element group 96:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_entry_sample_req_ps
      -- CP-element group 96: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_entry_sample_req
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:phi_stmt_1854_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1854_entry_sample_req_4897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1854_entry_sample_req_4897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(96), ack => phi_stmt_1854_req_0); -- 
    -- Element group maxPool3D_CP_4436_elements(96) is bound as output of CP function.
    -- CP-element group 97:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_phi_mux_ack_ps
      -- CP-element group 97: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/phi_stmt_1854_phi_mux_ack
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:phi_stmt_1854_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1854_phi_mux_ack_4900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1854_ack_0, ack => maxPool3D_CP_4436_elements(97)); -- 
    -- CP-element group 98:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (4) 
      -- CP-element group 98: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_chlx_x0_at_entry_1856_sample_completed__ps
      -- CP-element group 98: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_chlx_x0_at_entry_1856_sample_start__ps
      -- CP-element group 98: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_chlx_x0_at_entry_1856_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_chlx_x0_at_entry_1856_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(98) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_chlx_x0_at_entry_1856_update_start__ps
      -- CP-element group 99: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_chlx_x0_at_entry_1856_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(99) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(99) is bound as output of CP function.
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_chlx_x0_at_entry_1856_update_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(100) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(100) <= maxPool3D_CP_4436_elements(101);
    -- CP-element group 101:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	100 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/R_chlx_x0_at_entry_1856_update_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(101) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => maxPool3D_CP_4436_elements(99), ack => maxPool3D_CP_4436_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_sample_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(102) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_update_start__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(103) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_Sample/rr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1858_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(104), ack => type_cast_1858_inst_req_0); -- 
    maxPool3D_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(102) & maxPool3D_CP_4436_elements(106);
      gj_maxPool3D_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_update_start_
      -- CP-element group 105: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_Update/cr
      -- CP-element group 105: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_Update/$entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1858_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(105), ack => type_cast_1858_inst_req_1); -- 
    maxPool3D_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(103) & maxPool3D_CP_4436_elements(107);
      gj_maxPool3D_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	104 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_Sample/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1858_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1858_inst_ack_0, ack => maxPool3D_CP_4436_elements(106)); -- 
    -- CP-element group 107:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1858_update_completed__ps
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1858_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1858_inst_ack_1, ack => maxPool3D_CP_4436_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	92 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1862_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(108), ack => type_cast_1862_inst_req_0); -- 
    maxPool3D_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(92) & maxPool3D_CP_4436_elements(110);
      gj_maxPool3D_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	122 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_Update/cr
      -- CP-element group 109: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_Update/$entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1862_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(109), ack => type_cast_1862_inst_req_1); -- 
    maxPool3D_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(111) & maxPool3D_CP_4436_elements(122);
      gj_maxPool3D_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	88 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_Sample/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1862_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1862_inst_ack_0, ack => maxPool3D_CP_4436_elements(110)); -- 
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	120 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1862_Update/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1862_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1862_inst_ack_1, ack => maxPool3D_CP_4436_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	71 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1866_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(112), ack => type_cast_1866_inst_req_0); -- 
    maxPool3D_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(71) & maxPool3D_CP_4436_elements(114);
      gj_maxPool3D_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: 	122 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_Update/cr
      -- CP-element group 113: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1866_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(113), ack => type_cast_1866_inst_req_1); -- 
    maxPool3D_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(115) & maxPool3D_CP_4436_elements(122);
      gj_maxPool3D_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	67 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_sample_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1866_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1866_inst_ack_0, ack => maxPool3D_CP_4436_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	120 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1866_update_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1866_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1866_inst_ack_1, ack => maxPool3D_CP_4436_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	50 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1870_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(116), ack => type_cast_1870_inst_req_0); -- 
    maxPool3D_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(50) & maxPool3D_CP_4436_elements(118);
      gj_maxPool3D_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: 	122 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_Update/cr
      -- CP-element group 117: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1870_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(117), ack => type_cast_1870_inst_req_1); -- 
    maxPool3D_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(119) & maxPool3D_CP_4436_elements(122);
      gj_maxPool3D_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	48 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_Sample/ra
      -- CP-element group 118: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_sample_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(118) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1870_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1870_inst_ack_0, ack => maxPool3D_CP_4436_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	117 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_Update/ca
      -- CP-element group 119: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1870_update_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1870_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1870_inst_ack_1, ack => maxPool3D_CP_4436_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	111 
    -- CP-element group 120: 	115 
    -- CP-element group 120: 	119 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_Sample/crr
      -- CP-element group 120: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1939_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_4978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(120), ack => call_stmt_1939_call_req_0); -- 
    maxPool3D_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(111) & maxPool3D_CP_4436_elements(115) & maxPool3D_CP_4436_elements(119) & maxPool3D_CP_4436_elements(122);
      gj_maxPool3D_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_Update/ccr
      -- CP-element group 121: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1939_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_4983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(121), ack => call_stmt_1939_call_req_1); -- 
    maxPool3D_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool3D_CP_4436_elements(123);
      gj_maxPool3D_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	109 
    -- CP-element group 122: 	113 
    -- CP-element group 122: 	117 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_Sample/cra
      -- CP-element group 122: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_sample_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(122) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1939_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_4979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1939_call_ack_0, ack => maxPool3D_CP_4436_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	161 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	121 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_Update/cca
      -- CP-element group 123: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/call_stmt_1939_update_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_1939_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_4984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1939_call_ack_1, ack => maxPool3D_CP_4436_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	92 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_Sample/rr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1948_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(124), ack => type_cast_1948_inst_req_0); -- 
    maxPool3D_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(92) & maxPool3D_CP_4436_elements(126);
      gj_maxPool3D_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	44 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: 	130 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_update_start_
      -- CP-element group 125: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_Update/cr
      -- CP-element group 125: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_Update/$entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1948_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(125), ack => type_cast_1948_inst_req_1); -- 
    maxPool3D_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(44) & maxPool3D_CP_4436_elements(127) & maxPool3D_CP_4436_elements(130);
      gj_maxPool3D_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	88 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_Sample/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1948_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1948_inst_ack_0, ack => maxPool3D_CP_4436_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	87 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_Update/ca
      -- CP-element group 127: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1948_Update/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1948_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1948_inst_ack_1, ack => maxPool3D_CP_4436_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1957_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(128), ack => type_cast_1957_inst_req_0); -- 
    maxPool3D_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(127) & maxPool3D_CP_4436_elements(130);
      gj_maxPool3D_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: 	142 
    -- CP-element group 129: 	154 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_update_start_
      -- CP-element group 129: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_Update/cr
      -- CP-element group 129: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_Update/$entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1957_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_5011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(129), ack => type_cast_1957_inst_req_1); -- 
    maxPool3D_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(131) & maxPool3D_CP_4436_elements(142) & maxPool3D_CP_4436_elements(154);
      gj_maxPool3D_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	125 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_Sample/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1957_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_0, ack => maxPool3D_CP_4436_elements(130)); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	140 
    -- CP-element group 131: 	152 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1957_Update/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(131) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1957_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_1, ack => maxPool3D_CP_4436_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	71 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_Sample/req
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(132) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_colx_x1_1949_delayed_2_0_1959_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_5020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(132), ack => W_colx_x1_1949_delayed_2_0_1959_inst_req_0); -- 
    maxPool3D_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(71) & maxPool3D_CP_4436_elements(134);
      gj_maxPool3D_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: 	142 
    -- CP-element group 133: 	154 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_update_start_
      -- CP-element group 133: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_Update/req
      -- CP-element group 133: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_Update/$entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(133) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_colx_x1_1949_delayed_2_0_1959_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_5025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(133), ack => W_colx_x1_1949_delayed_2_0_1959_inst_req_1); -- 
    maxPool3D_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(135) & maxPool3D_CP_4436_elements(142) & maxPool3D_CP_4436_elements(154);
      gj_maxPool3D_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	67 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_Sample/ack
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(134) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_colx_x1_1949_delayed_2_0_1959_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1_1949_delayed_2_0_1959_inst_ack_0, ack => maxPool3D_CP_4436_elements(134)); -- 
    -- CP-element group 135:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	140 
    -- CP-element group 135: 	152 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_Update/ack
      -- CP-element group 135: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1961_Update/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(135) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_colx_x1_1949_delayed_2_0_1959_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1_1949_delayed_2_0_1959_inst_ack_1, ack => maxPool3D_CP_4436_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	92 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_Sample/req
      -- CP-element group 136: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(136) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_inc_1956_delayed_1_0_1967_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_5034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(136), ack => W_inc_1956_delayed_1_0_1967_inst_req_0); -- 
    maxPool3D_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(92) & maxPool3D_CP_4436_elements(138);
      gj_maxPool3D_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	44 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_Update/req
      -- CP-element group 137: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(137) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_inc_1956_delayed_1_0_1967_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_5039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(137), ack => W_inc_1956_delayed_1_0_1967_inst_req_1); -- 
    maxPool3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(44) & maxPool3D_CP_4436_elements(139);
      gj_maxPool3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	88 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_Sample/ack
      -- CP-element group 138: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_sample_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_inc_1956_delayed_1_0_1967_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inc_1956_delayed_1_0_1967_inst_ack_0, ack => maxPool3D_CP_4436_elements(138)); -- 
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	161 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	87 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_Update/ack
      -- CP-element group 139: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1969_update_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(139) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_inc_1956_delayed_1_0_1967_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inc_1956_delayed_1_0_1967_inst_ack_1, ack => maxPool3D_CP_4436_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	131 
    -- CP-element group 140: 	135 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_Sample/rr
      -- CP-element group 140: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1979_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(140), ack => type_cast_1979_inst_req_0); -- 
    maxPool3D_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(131) & maxPool3D_CP_4436_elements(135) & maxPool3D_CP_4436_elements(142);
      gj_maxPool3D_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	44 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: 	146 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_update_start_
      -- CP-element group 141: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_Update/$entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(141) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1979_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_5053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(141), ack => type_cast_1979_inst_req_1); -- 
    maxPool3D_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(44) & maxPool3D_CP_4436_elements(143) & maxPool3D_CP_4436_elements(146);
      gj_maxPool3D_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	129 
    -- CP-element group 142: 	133 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_Sample/ra
      -- CP-element group 142: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_Sample/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(142) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1979_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1979_inst_ack_0, ack => maxPool3D_CP_4436_elements(142)); -- 
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	66 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_Update/ca
      -- CP-element group 143: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1979_Update/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(143) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1979_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1979_inst_ack_1, ack => maxPool3D_CP_4436_elements(143)); -- 
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_Sample/rr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(144) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1988_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(144), ack => type_cast_1988_inst_req_0); -- 
    maxPool3D_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(143) & maxPool3D_CP_4436_elements(146);
      gj_maxPool3D_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	44 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: 	158 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_update_start_
      -- CP-element group 145: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_Update/cr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(145) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1988_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_5067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(145), ack => type_cast_1988_inst_req_1); -- 
    maxPool3D_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(44) & maxPool3D_CP_4436_elements(147) & maxPool3D_CP_4436_elements(158);
      gj_maxPool3D_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	141 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_Sample/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(146) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1988_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1988_inst_ack_0, ack => maxPool3D_CP_4436_elements(146)); -- 
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	156 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	47 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_1988_Update/ca
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(147) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_1988_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1988_inst_ack_1, ack => maxPool3D_CP_4436_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	50 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_Sample/req
      -- CP-element group 148: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_Sample/$entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(148) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_rowx_x1_1974_delayed_4_0_1990_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_5076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(148), ack => W_rowx_x1_1974_delayed_4_0_1990_inst_req_0); -- 
    maxPool3D_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(50) & maxPool3D_CP_4436_elements(150);
      gj_maxPool3D_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	44 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: 	158 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_Update/req
      -- CP-element group 149: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_update_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(149) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_rowx_x1_1974_delayed_4_0_1990_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_5081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(149), ack => W_rowx_x1_1974_delayed_4_0_1990_inst_req_1); -- 
    maxPool3D_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(44) & maxPool3D_CP_4436_elements(151) & maxPool3D_CP_4436_elements(158);
      gj_maxPool3D_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	48 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_Sample/ack
      -- CP-element group 150: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_sample_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(150) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_rowx_x1_1974_delayed_4_0_1990_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rowx_x1_1974_delayed_4_0_1990_inst_ack_0, ack => maxPool3D_CP_4436_elements(150)); -- 
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	156 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	47 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_Update/ack
      -- CP-element group 151: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_1992_Update/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(151) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_rowx_x1_1974_delayed_4_0_1990_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rowx_x1_1974_delayed_4_0_1990_inst_ack_1, ack => maxPool3D_CP_4436_elements(151)); -- 
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	131 
    -- CP-element group 152: 	135 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_Sample/req
      -- CP-element group 152: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_sample_start_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(152) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_5090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(152), ack => W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_req_0); -- 
    maxPool3D_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(131) & maxPool3D_CP_4436_elements(135) & maxPool3D_CP_4436_elements(154);
      gj_maxPool3D_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	44 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_update_start_
      -- CP-element group 153: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_Update/req
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(153) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_5095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(153), ack => W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_req_1); -- 
    maxPool3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(44) & maxPool3D_CP_4436_elements(155);
      gj_maxPool3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	129 
    -- CP-element group 154: 	133 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_Sample/ack
      -- CP-element group 154: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_sample_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(154) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_ack_0, ack => maxPool3D_CP_4436_elements(154)); -- 
    -- CP-element group 155:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	161 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	66 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/assign_stmt_2000_Update/ack
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(155) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_ack_1, ack => maxPool3D_CP_4436_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	147 
    -- CP-element group 156: 	151 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_Sample/rr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2010_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(156), ack => type_cast_2010_inst_req_0); -- 
    maxPool3D_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(147) & maxPool3D_CP_4436_elements(151) & maxPool3D_CP_4436_elements(158);
      gj_maxPool3D_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_update_start_
      -- CP-element group 157: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_Update/$entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2010_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_5109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(157), ack => type_cast_2010_inst_req_1); -- 
    maxPool3D_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool3D_CP_4436_elements(159);
      gj_maxPool3D_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	145 
    -- CP-element group 158: 	149 
    -- CP-element group 158: 	156 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_Sample/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(158) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2010_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2010_inst_ack_0, ack => maxPool3D_CP_4436_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	42 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/type_cast_2010_update_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2010_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2010_inst_ack_1, ack => maxPool3D_CP_4436_elements(159)); -- 
    -- CP-element group 160:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	41 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	42 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(160) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool3D_CP_4436_elements(160) is a control-delay.
    cp_element_160_delay: control_delay_element  generic map(name => " 160_delay", delay_value => 1)  port map(req => maxPool3D_CP_4436_elements(41), ack => maxPool3D_CP_4436_elements(160), clk => clk, reset =>reset);
    -- CP-element group 161:  join  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	123 
    -- CP-element group 161: 	139 
    -- CP-element group 161: 	155 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	38 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1711/do_while_stmt_1842/do_while_stmt_1842_loop_body/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(161) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_4436_elements(123) & maxPool3D_CP_4436_elements(139) & maxPool3D_CP_4436_elements(155);
      gj_maxPool3D_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_4436_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	37 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_1711/do_while_stmt_1842/loop_exit/ack
      -- CP-element group 162: 	 branch_block_stmt_1711/do_while_stmt_1842/loop_exit/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:do_while_stmt_1842_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1842_branch_ack_0, ack => maxPool3D_CP_4436_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	37 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_1711/do_while_stmt_1842/loop_taken/$exit
      -- CP-element group 163: 	 branch_block_stmt_1711/do_while_stmt_1842/loop_taken/ack
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:do_while_stmt_1842_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1842_branch_ack_1, ack => maxPool3D_CP_4436_elements(163)); -- 
    -- CP-element group 164:  transition  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	35 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	1 
    -- CP-element group 164:  members (1) 
      -- CP-element group 164: 	 branch_block_stmt_1711/do_while_stmt_1842/$exit
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(164) fired."); 
        -- 
      end if; --
    end process; 
    maxPool3D_CP_4436_elements(164) <= maxPool3D_CP_4436_elements(35);
    -- CP-element group 165:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	1 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: 	168 
    -- CP-element group 165:  members (18) 
      -- CP-element group 165: 	 branch_block_stmt_1711/assign_stmt_2032__entry__
      -- CP-element group 165: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_Update/cr
      -- CP-element group 165: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_Update/$entry
      -- CP-element group 165: 	 branch_block_stmt_1711/assign_stmt_2032/$entry
      -- CP-element group 165: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_Sample/rr
      -- CP-element group 165: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_1711/merge_stmt_2027__exit__
      -- CP-element group 165: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_update_start_
      -- CP-element group 165: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_1711/if_stmt_2023_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_1711/if_stmt_2023_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_1711/whilex_xbody_whilex_xend
      -- CP-element group 165: 	 branch_block_stmt_1711/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_1711/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_1711/merge_stmt_2027_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_1711/merge_stmt_2027_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_1711/merge_stmt_2027_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_1711/merge_stmt_2027_PhiAck/dummy
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:if_stmt_2023_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2031_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2031_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_5133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2023_branch_ack_1, ack => maxPool3D_CP_4436_elements(165)); -- 
    cr_5154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(165), ack => type_cast_2031_inst_req_1); -- 
    rr_5149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(165), ack => type_cast_2031_inst_req_0); -- 
    -- CP-element group 166:  merge  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	1 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (5) 
      -- CP-element group 166: 	 branch_block_stmt_1711/if_stmt_2023__exit__
      -- CP-element group 166: 	 branch_block_stmt_1711/merge_stmt_2027__entry__
      -- CP-element group 166: 	 branch_block_stmt_1711/if_stmt_2023_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_1711/if_stmt_2023_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_1711/merge_stmt_2027_dead_link/$entry
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(166) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:if_stmt_2023_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_5137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2023_branch_ack_0, ack => maxPool3D_CP_4436_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_sample_completed_
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2031_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2031_inst_ack_0, ack => maxPool3D_CP_4436_elements(167)); -- 
    -- CP-element group 168:  fork  transition  place  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	165 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168: 	170 
    -- CP-element group 168: 	172 
    -- CP-element group 168:  members (16) 
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048__entry__
      -- CP-element group 168: 	 branch_block_stmt_1711/assign_stmt_2032/$exit
      -- CP-element group 168: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_1711/assign_stmt_2032__exit__
      -- CP-element group 168: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_1711/assign_stmt_2032/type_cast_2031_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_update_start_
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/$entry
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_Sample/crr
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_Update/ccr
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_update_start_
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_Update/cr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(168)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(168)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(168) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2031_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_2035_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_2035_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2039_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2031_inst_ack_1, ack => maxPool3D_CP_4436_elements(168)); -- 
    crr_5166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(168), ack => call_stmt_2035_call_req_0); -- 
    ccr_5171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(168), ack => call_stmt_2035_call_req_1); -- 
    cr_5185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(168), ack => type_cast_2039_inst_req_1); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_Sample/cra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(169)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(169)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(169) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_2035_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_5167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2035_call_ack_0, ack => maxPool3D_CP_4436_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (6) 
      -- CP-element group 170: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/call_stmt_2035_Update/cca
      -- CP-element group 170: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_Sample/rr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(170)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(170)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(170) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_2035_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2039_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_5172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2035_call_ack_1, ack => maxPool3D_CP_4436_elements(170)); -- 
    rr_5180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(170), ack => type_cast_2039_inst_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_Sample/ra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(171)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(171)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(171) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2039_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2039_inst_ack_0, ack => maxPool3D_CP_4436_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	168 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (6) 
      -- CP-element group 172: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/type_cast_2039_Update/ca
      -- CP-element group 172: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_Sample/req
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(172)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(172)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(172) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:type_cast_2039_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:WPIPE_elapsed_time_pipe_2046_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_5186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2039_inst_ack_1, ack => maxPool3D_CP_4436_elements(172)); -- 
    req_5194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(172), ack => WPIPE_elapsed_time_pipe_2046_inst_req_0); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_update_start_
      -- CP-element group 173: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_Sample/ack
      -- CP-element group 173: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_Update/req
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(173)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(173)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(173) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:WPIPE_elapsed_time_pipe_2046_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:WPIPE_elapsed_time_pipe_2046_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_2046_inst_ack_0, ack => maxPool3D_CP_4436_elements(173)); -- 
    req_5199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(173), ack => WPIPE_elapsed_time_pipe_2046_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  place  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (13) 
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048__exit__
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2050__entry__
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/$exit
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2035_to_assign_stmt_2048/WPIPE_elapsed_time_pipe_2046_Update/ack
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2050/$entry
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_update_start_
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_Sample/crr
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_Update/ccr
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(174)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(174)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(174) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:WPIPE_elapsed_time_pipe_2046_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_2050_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_2050_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_2046_inst_ack_1, ack => maxPool3D_CP_4436_elements(174)); -- 
    crr_5211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(174), ack => call_stmt_2050_call_req_0); -- 
    ccr_5216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_4436_elements(174), ack => call_stmt_2050_call_req_1); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_Sample/cra
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(175)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(175)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(175) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_2050_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_5212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2050_call_ack_0, ack => maxPool3D_CP_4436_elements(175)); -- 
    -- CP-element group 176:  transition  place  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (16) 
      -- CP-element group 176: 	 branch_block_stmt_1711/return__
      -- CP-element group 176: 	 branch_block_stmt_1711/merge_stmt_2052__exit__
      -- CP-element group 176: 	 branch_block_stmt_1711/call_stmt_2050__exit__
      -- CP-element group 176: 	 branch_block_stmt_1711/branch_block_stmt_1711__exit__
      -- CP-element group 176: 	 $exit
      -- CP-element group 176: 	 branch_block_stmt_1711/$exit
      -- CP-element group 176: 	 branch_block_stmt_1711/call_stmt_2050/$exit
      -- CP-element group 176: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_1711/call_stmt_2050/call_stmt_2050_Update/cca
      -- CP-element group 176: 	 branch_block_stmt_1711/return___PhiReq/$entry
      -- CP-element group 176: 	 branch_block_stmt_1711/return___PhiReq/$exit
      -- CP-element group 176: 	 branch_block_stmt_1711/merge_stmt_2052_PhiReqMerge
      -- CP-element group 176: 	 branch_block_stmt_1711/merge_stmt_2052_PhiAck/$entry
      -- CP-element group 176: 	 branch_block_stmt_1711/merge_stmt_2052_PhiAck/$exit
      -- CP-element group 176: 	 branch_block_stmt_1711/merge_stmt_2052_PhiAck/dummy
      -- 
    -- logger for CP element group maxPool3D_CP_4436_elements(176)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool3D_CP_4436_elements(176)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:maxPool3D_CP_4436_elements(176) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool3D:CP:call_stmt_2050_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_5217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2050_call_ack_1, ack => maxPool3D_CP_4436_elements(176)); -- 
    maxPool3D_do_while_stmt_1842_terminator_5120: loop_terminator -- 
      generic map (name => " maxPool3D_do_while_stmt_1842_terminator_5120", max_iterations_in_flight =>15) 
      port map(loop_body_exit => maxPool3D_CP_4436_elements(38),loop_continue => maxPool3D_CP_4436_elements(163),loop_terminate => maxPool3D_CP_4436_elements(162),loop_back => maxPool3D_CP_4436_elements(36),loop_exit => maxPool3D_CP_4436_elements(35),clk => clk, reset => reset); -- 
    phi_stmt_1844_phi_seq_4840_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_4436_elements(51);
      maxPool3D_CP_4436_elements(56)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_4436_elements(60);
      maxPool3D_CP_4436_elements(57)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_4436_elements(61);
      maxPool3D_CP_4436_elements(52) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_4436_elements(53);
      maxPool3D_CP_4436_elements(62)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_4436_elements(62);
      maxPool3D_CP_4436_elements(63)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_4436_elements(64);
      maxPool3D_CP_4436_elements(54) <= phi_mux_reqs(1);
      phi_stmt_1844_phi_seq_4840 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1844_phi_seq_4840") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_4436_elements(43), 
          phi_sample_ack => maxPool3D_CP_4436_elements(49), 
          phi_update_req => maxPool3D_CP_4436_elements(45), 
          phi_update_ack => maxPool3D_CP_4436_elements(50), 
          phi_mux_ack => maxPool3D_CP_4436_elements(55), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1849_phi_seq_4884_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_4436_elements(72);
      maxPool3D_CP_4436_elements(77)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_4436_elements(81);
      maxPool3D_CP_4436_elements(78)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_4436_elements(82);
      maxPool3D_CP_4436_elements(73) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_4436_elements(74);
      maxPool3D_CP_4436_elements(83)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_4436_elements(83);
      maxPool3D_CP_4436_elements(84)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_4436_elements(85);
      maxPool3D_CP_4436_elements(75) <= phi_mux_reqs(1);
      phi_stmt_1849_phi_seq_4884 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1849_phi_seq_4884") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_4436_elements(68), 
          phi_sample_ack => maxPool3D_CP_4436_elements(69), 
          phi_update_req => maxPool3D_CP_4436_elements(70), 
          phi_update_ack => maxPool3D_CP_4436_elements(71), 
          phi_mux_ack => maxPool3D_CP_4436_elements(76), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1854_phi_seq_4928_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_4436_elements(95);
      maxPool3D_CP_4436_elements(98)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_4436_elements(98);
      maxPool3D_CP_4436_elements(99)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_4436_elements(100);
      maxPool3D_CP_4436_elements(96) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_4436_elements(93);
      maxPool3D_CP_4436_elements(102)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_4436_elements(106);
      maxPool3D_CP_4436_elements(103)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_4436_elements(107);
      maxPool3D_CP_4436_elements(94) <= phi_mux_reqs(1);
      phi_stmt_1854_phi_seq_4928 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1854_phi_seq_4928") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_4436_elements(89), 
          phi_sample_ack => maxPool3D_CP_4436_elements(90), 
          phi_update_req => maxPool3D_CP_4436_elements(91), 
          phi_update_ack => maxPool3D_CP_4436_elements(92), 
          phi_mux_ack => maxPool3D_CP_4436_elements(97), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4792_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= maxPool3D_CP_4436_elements(39);
        preds(1)  <= maxPool3D_CP_4436_elements(40);
        entry_tmerge_4792 : transition_merge -- 
          generic map(name => " entry_tmerge_4792")
          port map (preds => preds, symbol_out => maxPool3D_CP_4436_elements(41));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_2022_wire : std_logic_vector(0 downto 0);
    signal add43_1881 : std_logic_vector(31 downto 0);
    signal add45_1891 : std_logic_vector(31 downto 0);
    signal add57_1907 : std_logic_vector(31 downto 0);
    signal add60_1917 : std_logic_vector(31 downto 0);
    signal add67_1922 : std_logic_vector(31 downto 0);
    signal add71_1927 : std_logic_vector(31 downto 0);
    signal add74_1932 : std_logic_vector(31 downto 0);
    signal add_1817 : std_logic_vector(31 downto 0);
    signal call103_2035 : std_logic_vector(63 downto 0);
    signal call75_1939 : std_logic_vector(7 downto 0);
    signal call_1787 : std_logic_vector(63 downto 0);
    signal chlx_x0_1854 : std_logic_vector(15 downto 0);
    signal chlx_x0_at_entry_1836 : std_logic_vector(15 downto 0);
    signal chlx_x1_1976 : std_logic_vector(15 downto 0);
    signal cmp88_1985 : std_logic_vector(0 downto 0);
    signal cmp98_2016 : std_logic_vector(0 downto 0);
    signal cmp_1954 : std_logic_vector(0 downto 0);
    signal colx_x1_1849 : std_logic_vector(15 downto 0);
    signal colx_x1_1949_delayed_2_0_1961 : std_logic_vector(15 downto 0);
    signal colx_x1_at_entry_1831 : std_logic_vector(15 downto 0);
    signal colx_x2_2007 : std_logic_vector(15 downto 0);
    signal conv104_2040 : std_logic_vector(63 downto 0);
    signal conv12_1773 : std_logic_vector(31 downto 0);
    signal conv14_1779 : std_logic_vector(31 downto 0);
    signal conv17_2032 : std_logic_vector(63 downto 0);
    signal conv27_1794 : std_logic_vector(31 downto 0);
    signal conv33_1863 : std_logic_vector(31 downto 0);
    signal conv37_1867 : std_logic_vector(31 downto 0);
    signal conv39_1800 : std_logic_vector(31 downto 0);
    signal conv41_1871 : std_logic_vector(31 downto 0);
    signal conv78_1949 : std_logic_vector(31 downto 0);
    signal conv85_1980 : std_logic_vector(31 downto 0);
    signal conv95_2011 : std_logic_vector(31 downto 0);
    signal conv97_1823 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1721 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1733 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1745 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1757 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1806 : std_logic_vector(31 downto 0);
    signal inc83_1958 : std_logic_vector(15 downto 0);
    signal inc83x_xcolx_x1_1966 : std_logic_vector(15 downto 0);
    signal inc83x_xcolx_x1_1981_delayed_1_0_2000 : std_logic_vector(15 downto 0);
    signal inc92_1989 : std_logic_vector(15 downto 0);
    signal inc92x_xrowx_x1_1997 : std_logic_vector(15 downto 0);
    signal inc_1945 : std_logic_vector(15 downto 0);
    signal inc_1956_delayed_1_0_1969 : std_logic_vector(15 downto 0);
    signal mul42_1876 : std_logic_vector(31 downto 0);
    signal mul44_1886 : std_logic_vector(31 downto 0);
    signal mul56_1902 : std_logic_vector(31 downto 0);
    signal mul58_1812 : std_logic_vector(31 downto 0);
    signal mul_1784 : std_logic_vector(31 downto 0);
    signal ptr_deref_1724_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1724_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1724_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1724_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1724_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1736_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1736_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1736_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1736_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1736_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1748_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1748_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1748_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1748_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1748_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1748_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1748_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1748_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_1748_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_1748_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_1748_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1748_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_1748_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_1748_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_1760_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1760_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1760_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1760_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1760_word_offset_0 : std_logic_vector(6 downto 0);
    signal rowx_x1_1844 : std_logic_vector(15 downto 0);
    signal rowx_x1_1974_delayed_4_0_1992 : std_logic_vector(15 downto 0);
    signal rowx_x1_at_entry_1826 : std_logic_vector(15 downto 0);
    signal shl59_1912 : std_logic_vector(31 downto 0);
    signal shl_1897 : std_logic_vector(31 downto 0);
    signal shr_1767 : std_logic_vector(31 downto 0);
    signal sub_2045 : std_logic_vector(63 downto 0);
    signal tmp2_1737 : std_logic_vector(31 downto 0);
    signal tmp5_1749 : std_logic_vector(31 downto 0);
    signal tmp8_1761 : std_logic_vector(31 downto 0);
    signal tmp_1725 : std_logic_vector(31 downto 0);
    signal type_cast_1765_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1771_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1777_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1792_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1798_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1804_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1810_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1821_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1847_wire : std_logic_vector(15 downto 0);
    signal type_cast_1852_wire : std_logic_vector(15 downto 0);
    signal type_cast_1858_wire : std_logic_vector(15 downto 0);
    signal type_cast_1895_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1943_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1973_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2004_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2030_wire : std_logic_vector(63 downto 0);
    signal type_cast_2038_wire : std_logic_vector(63 downto 0);
    signal whilex_xbody_whilex_xend_taken_2019 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    chlx_x0_at_entry_1836 <= "0000000000000000";
    colx_x1_at_entry_1831 <= "0000000000000000";
    iNsTr_2_1721 <= "00000000000000000000000000000011";
    iNsTr_3_1733 <= "00000000000000000000000000000010";
    iNsTr_4_1745 <= "00000000000000000000000000001101";
    iNsTr_5_1757 <= "00000000000000000000000000000100";
    ptr_deref_1724_word_offset_0 <= "0000000";
    ptr_deref_1736_word_offset_0 <= "0000000";
    ptr_deref_1748_word_offset_0 <= "000000000";
    ptr_deref_1748_word_offset_1 <= "000000001";
    ptr_deref_1748_word_offset_2 <= "000000010";
    ptr_deref_1748_word_offset_3 <= "000000011";
    ptr_deref_1760_word_offset_0 <= "0000000";
    rowx_x1_at_entry_1826 <= "0000000000000000";
    type_cast_1765_wire_constant <= "00000000000000000000000000000100";
    type_cast_1771_wire_constant <= "00000000000000001111111111111111";
    type_cast_1777_wire_constant <= "00000000000000001111111111111111";
    type_cast_1792_wire_constant <= "00000000000000001111111111111111";
    type_cast_1798_wire_constant <= "00000000000000001111111111111111";
    type_cast_1804_wire_constant <= "00000000000000000000000000000011";
    type_cast_1810_wire_constant <= "00000000000000011111111111111110";
    type_cast_1821_wire_constant <= "00000000000000001111111111111111";
    type_cast_1895_wire_constant <= "00000000000000000000000000000010";
    type_cast_1943_wire_constant <= "0000000000000001";
    type_cast_1973_wire_constant <= "0000000000000000";
    type_cast_2004_wire_constant <= "0000000000000000";
    -- logger for phi phi_stmt_1844
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1844_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:maxPool3D:DP:phi_stmt_1844:input-0 type_cast_1847_wire= " & Convert_SLV_To_Hex_String(type_cast_1847_wire));
          --
        end if;
        if phi_stmt_1844_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:maxPool3D:DP:phi_stmt_1844:input-1 rowx_x1_at_entry_1826= " & Convert_SLV_To_Hex_String(rowx_x1_at_entry_1826));
          --
        end if;
        if phi_stmt_1844_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:maxPool3D:DP:phi_stmt_1844:sample-completed");
          --
        end if;
        if phi_stmt_1844_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:maxPool3D:DP:phi_stmt_1844:output rowx_x1_1844= " & Convert_SLV_To_Hex_String(rowx_x1_1844));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1844: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1847_wire & rowx_x1_at_entry_1826;
      req <= phi_stmt_1844_req_0 & phi_stmt_1844_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1844",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1844_ack_0,
          idata => idata,
          odata => rowx_x1_1844,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1844
    -- logger for phi phi_stmt_1849
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1849_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:maxPool3D:DP:phi_stmt_1849:input-0 type_cast_1852_wire= " & Convert_SLV_To_Hex_String(type_cast_1852_wire));
          --
        end if;
        if phi_stmt_1849_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:maxPool3D:DP:phi_stmt_1849:input-1 colx_x1_at_entry_1831= " & Convert_SLV_To_Hex_String(colx_x1_at_entry_1831));
          --
        end if;
        if phi_stmt_1849_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:maxPool3D:DP:phi_stmt_1849:sample-completed");
          --
        end if;
        if phi_stmt_1849_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:maxPool3D:DP:phi_stmt_1849:output colx_x1_1849= " & Convert_SLV_To_Hex_String(colx_x1_1849));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1849: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1852_wire & colx_x1_at_entry_1831;
      req <= phi_stmt_1849_req_0 & phi_stmt_1849_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1849",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1849_ack_0,
          idata => idata,
          odata => colx_x1_1849,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1849
    -- logger for phi phi_stmt_1854
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1854_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:maxPool3D:DP:phi_stmt_1854:input-0 chlx_x0_at_entry_1836= " & Convert_SLV_To_Hex_String(chlx_x0_at_entry_1836));
          --
        end if;
        if phi_stmt_1854_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:maxPool3D:DP:phi_stmt_1854:input-1 type_cast_1858_wire= " & Convert_SLV_To_Hex_String(type_cast_1858_wire));
          --
        end if;
        if phi_stmt_1854_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:maxPool3D:DP:phi_stmt_1854:sample-completed");
          --
        end if;
        if phi_stmt_1854_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:maxPool3D:DP:phi_stmt_1854:output chlx_x0_1854= " & Convert_SLV_To_Hex_String(chlx_x0_1854));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1854: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= chlx_x0_at_entry_1836 & type_cast_1858_wire;
      req <= phi_stmt_1854_req_0 & phi_stmt_1854_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1854",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1854_ack_0,
          idata => idata,
          odata => chlx_x0_1854,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1854
    -- logger for split-operator MUX_1975_inst flow-through 
    process(chlx_x1_1976) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:MUX_1975_inst:flowthrough inputs: " & " cmp_1954 = "& Convert_SLV_To_Hex_String(cmp_1954) & " type_cast_1973_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1973_wire_constant) & " inc_1956_delayed_1_0_1969 = "& Convert_SLV_To_Hex_String(inc_1956_delayed_1_0_1969) & " outputs:" & " chlx_x1_1976= "  & Convert_SLV_To_Hex_String(chlx_x1_1976));
      --
    end process; 
    -- flow-through select operator MUX_1975_inst
    chlx_x1_1976 <= type_cast_1973_wire_constant when (cmp_1954(0) /=  '0') else inc_1956_delayed_1_0_1969;
    -- logger for split-operator MUX_2006_inst flow-through 
    process(colx_x2_2007) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:MUX_2006_inst:flowthrough inputs: " & " cmp88_1985 = "& Convert_SLV_To_Hex_String(cmp88_1985) & " type_cast_2004_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_2004_wire_constant) & " inc83x_xcolx_x1_1981_delayed_1_0_2000 = "& Convert_SLV_To_Hex_String(inc83x_xcolx_x1_1981_delayed_1_0_2000) & " outputs:" & " colx_x2_2007= "  & Convert_SLV_To_Hex_String(colx_x2_2007));
      --
    end process; 
    -- flow-through select operator MUX_2006_inst
    colx_x2_2007 <= type_cast_2004_wire_constant when (cmp88_1985(0) /=  '0') else inc83x_xcolx_x1_1981_delayed_1_0_2000;
    -- logger for split-operator W_colx_x1_1949_delayed_2_0_1959_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_colx_x1_1949_delayed_2_0_1959_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:W_colx_x1_1949_delayed_2_0_1959_inst:started:   inputs: " & " colx_x1_1849 = "& Convert_SLV_To_Hex_String(colx_x1_1849));
          --
        end if; 
        if W_colx_x1_1949_delayed_2_0_1959_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:W_colx_x1_1949_delayed_2_0_1959_inst:finished:  outputs: " & " colx_x1_1949_delayed_2_0_1961= "  & Convert_SLV_To_Hex_String(colx_x1_1949_delayed_2_0_1961));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_colx_x1_1949_delayed_2_0_1959_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_colx_x1_1949_delayed_2_0_1959_inst_req_0;
      W_colx_x1_1949_delayed_2_0_1959_inst_ack_0<= wack(0);
      rreq(0) <= W_colx_x1_1949_delayed_2_0_1959_inst_req_1;
      W_colx_x1_1949_delayed_2_0_1959_inst_ack_1<= rack(0);
      W_colx_x1_1949_delayed_2_0_1959_inst : InterlockBuffer generic map ( -- 
        name => "W_colx_x1_1949_delayed_2_0_1959_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1_1849,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => colx_x1_1949_delayed_2_0_1961,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst:started:   inputs: " & " inc83x_xcolx_x1_1966 = "& Convert_SLV_To_Hex_String(inc83x_xcolx_x1_1966));
          --
        end if; 
        if W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst:finished:  outputs: " & " inc83x_xcolx_x1_1981_delayed_1_0_2000= "  & Convert_SLV_To_Hex_String(inc83x_xcolx_x1_1981_delayed_1_0_2000));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_req_0;
      W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_ack_0<= wack(0);
      rreq(0) <= W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_req_1;
      W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst_ack_1<= rack(0);
      W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst : InterlockBuffer generic map ( -- 
        name => "W_inc83x_xcolx_x1_1981_delayed_1_0_1998_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc83x_xcolx_x1_1966,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc83x_xcolx_x1_1981_delayed_1_0_2000,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_inc_1956_delayed_1_0_1967_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_inc_1956_delayed_1_0_1967_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:W_inc_1956_delayed_1_0_1967_inst:started:   inputs: " & " inc_1945 = "& Convert_SLV_To_Hex_String(inc_1945));
          --
        end if; 
        if W_inc_1956_delayed_1_0_1967_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:W_inc_1956_delayed_1_0_1967_inst:finished:  outputs: " & " inc_1956_delayed_1_0_1969= "  & Convert_SLV_To_Hex_String(inc_1956_delayed_1_0_1969));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_inc_1956_delayed_1_0_1967_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_inc_1956_delayed_1_0_1967_inst_req_0;
      W_inc_1956_delayed_1_0_1967_inst_ack_0<= wack(0);
      rreq(0) <= W_inc_1956_delayed_1_0_1967_inst_req_1;
      W_inc_1956_delayed_1_0_1967_inst_ack_1<= rack(0);
      W_inc_1956_delayed_1_0_1967_inst : InterlockBuffer generic map ( -- 
        name => "W_inc_1956_delayed_1_0_1967_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_1945,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_1956_delayed_1_0_1969,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_rowx_x1_1974_delayed_4_0_1990_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_rowx_x1_1974_delayed_4_0_1990_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:W_rowx_x1_1974_delayed_4_0_1990_inst:started:   inputs: " & " rowx_x1_1844 = "& Convert_SLV_To_Hex_String(rowx_x1_1844));
          --
        end if; 
        if W_rowx_x1_1974_delayed_4_0_1990_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:W_rowx_x1_1974_delayed_4_0_1990_inst:finished:  outputs: " & " rowx_x1_1974_delayed_4_0_1992= "  & Convert_SLV_To_Hex_String(rowx_x1_1974_delayed_4_0_1992));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_rowx_x1_1974_delayed_4_0_1990_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rowx_x1_1974_delayed_4_0_1990_inst_req_0;
      W_rowx_x1_1974_delayed_4_0_1990_inst_ack_0<= wack(0);
      rreq(0) <= W_rowx_x1_1974_delayed_4_0_1990_inst_req_1;
      W_rowx_x1_1974_delayed_4_0_1990_inst_ack_1<= rack(0);
      W_rowx_x1_1974_delayed_4_0_1990_inst : InterlockBuffer generic map ( -- 
        name => "W_rowx_x1_1974_delayed_4_0_1990_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rowx_x1_1844,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rowx_x1_1974_delayed_4_0_1992,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_whilex_xbody_whilex_xend_taken_2017_inst flow-through 
    process(whilex_xbody_whilex_xend_taken_2019) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:W_whilex_xbody_whilex_xend_taken_2017_inst:flowthrough inputs: " & " cmp98_2016 = "& Convert_SLV_To_Hex_String(cmp98_2016) & " outputs:" & " whilex_xbody_whilex_xend_taken_2019= "  & Convert_SLV_To_Hex_String(whilex_xbody_whilex_xend_taken_2019));
      --
    end process; 
    -- interlock W_whilex_xbody_whilex_xend_taken_2017_inst
    process(cmp98_2016) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp98_2016(0 downto 0);
      whilex_xbody_whilex_xend_taken_2019 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1847_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1847_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1847_inst:started:   inputs: " & " inc92x_xrowx_x1_1997 = "& Convert_SLV_To_Hex_String(inc92x_xrowx_x1_1997));
          --
        end if; 
        if type_cast_1847_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1847_inst:finished:  outputs: " & " type_cast_1847_wire= "  & Convert_SLV_To_Hex_String(type_cast_1847_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1847_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1847_inst_req_0;
      type_cast_1847_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1847_inst_req_1;
      type_cast_1847_inst_ack_1<= rack(0);
      type_cast_1847_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1847_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc92x_xrowx_x1_1997,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1847_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1852_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1852_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1852_inst:started:   inputs: " & " colx_x2_2007 = "& Convert_SLV_To_Hex_String(colx_x2_2007));
          --
        end if; 
        if type_cast_1852_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1852_inst:finished:  outputs: " & " type_cast_1852_wire= "  & Convert_SLV_To_Hex_String(type_cast_1852_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1852_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1852_inst_req_0;
      type_cast_1852_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1852_inst_req_1;
      type_cast_1852_inst_ack_1<= rack(0);
      type_cast_1852_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1852_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x2_2007,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1852_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1858_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1858_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1858_inst:started:   inputs: " & " chlx_x1_1976 = "& Convert_SLV_To_Hex_String(chlx_x1_1976));
          --
        end if; 
        if type_cast_1858_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1858_inst:finished:  outputs: " & " type_cast_1858_wire= "  & Convert_SLV_To_Hex_String(type_cast_1858_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1858_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1858_inst_req_0;
      type_cast_1858_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1858_inst_req_1;
      type_cast_1858_inst_ack_1<= rack(0);
      type_cast_1858_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1858_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x1_1976,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1858_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1862_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1862_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1862_inst:started:   inputs: " & " chlx_x0_1854 = "& Convert_SLV_To_Hex_String(chlx_x0_1854));
          --
        end if; 
        if type_cast_1862_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1862_inst:finished:  outputs: " & " conv33_1863= "  & Convert_SLV_To_Hex_String(conv33_1863));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1862_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1862_inst_req_0;
      type_cast_1862_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1862_inst_req_1;
      type_cast_1862_inst_ack_1<= rack(0);
      type_cast_1862_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1862_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x0_1854,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_1863,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1866_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1866_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1866_inst:started:   inputs: " & " colx_x1_1849 = "& Convert_SLV_To_Hex_String(colx_x1_1849));
          --
        end if; 
        if type_cast_1866_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1866_inst:finished:  outputs: " & " conv37_1867= "  & Convert_SLV_To_Hex_String(conv37_1867));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1866_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1866_inst_req_0;
      type_cast_1866_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1866_inst_req_1;
      type_cast_1866_inst_ack_1<= rack(0);
      type_cast_1866_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1866_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1_1849,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_1867,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1870_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1870_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1870_inst:started:   inputs: " & " rowx_x1_1844 = "& Convert_SLV_To_Hex_String(rowx_x1_1844));
          --
        end if; 
        if type_cast_1870_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1870_inst:finished:  outputs: " & " conv41_1871= "  & Convert_SLV_To_Hex_String(conv41_1871));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1870_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1870_inst_req_0;
      type_cast_1870_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1870_inst_req_1;
      type_cast_1870_inst_ack_1<= rack(0);
      type_cast_1870_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1870_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rowx_x1_1844,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_1871,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1948_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1948_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1948_inst:started:   inputs: " & " inc_1945 = "& Convert_SLV_To_Hex_String(inc_1945));
          --
        end if; 
        if type_cast_1948_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1948_inst:finished:  outputs: " & " conv78_1949= "  & Convert_SLV_To_Hex_String(conv78_1949));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1948_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1948_inst_req_0;
      type_cast_1948_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1948_inst_req_1;
      type_cast_1948_inst_ack_1<= rack(0);
      type_cast_1948_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1948_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_1945,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_1949,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1957_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1957_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1957_inst:started:   inputs: " & " cmp_1954 = "& Convert_SLV_To_Hex_String(cmp_1954));
          --
        end if; 
        if type_cast_1957_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1957_inst:finished:  outputs: " & " inc83_1958= "  & Convert_SLV_To_Hex_String(inc83_1958));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1957_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1957_inst_req_0;
      type_cast_1957_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1957_inst_req_1;
      type_cast_1957_inst_ack_1<= rack(0);
      type_cast_1957_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1957_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp_1954,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc83_1958,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1979_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1979_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1979_inst:started:   inputs: " & " inc83x_xcolx_x1_1966 = "& Convert_SLV_To_Hex_String(inc83x_xcolx_x1_1966));
          --
        end if; 
        if type_cast_1979_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1979_inst:finished:  outputs: " & " conv85_1980= "  & Convert_SLV_To_Hex_String(conv85_1980));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1979_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1979_inst_req_0;
      type_cast_1979_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1979_inst_req_1;
      type_cast_1979_inst_ack_1<= rack(0);
      type_cast_1979_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1979_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc83x_xcolx_x1_1966,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1980,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1988_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1988_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1988_inst:started:   inputs: " & " cmp88_1985 = "& Convert_SLV_To_Hex_String(cmp88_1985));
          --
        end if; 
        if type_cast_1988_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_1988_inst:finished:  outputs: " & " inc92_1989= "  & Convert_SLV_To_Hex_String(inc92_1989));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1988_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1988_inst_req_0;
      type_cast_1988_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1988_inst_req_1;
      type_cast_1988_inst_ack_1<= rack(0);
      type_cast_1988_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1988_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp88_1985,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc92_1989,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_2010_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_2010_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_2010_inst:started:   inputs: " & " inc92x_xrowx_x1_1997 = "& Convert_SLV_To_Hex_String(inc92x_xrowx_x1_1997));
          --
        end if; 
        if type_cast_2010_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_2010_inst:finished:  outputs: " & " conv95_2011= "  & Convert_SLV_To_Hex_String(conv95_2011));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_2010_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2010_inst_req_0;
      type_cast_2010_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2010_inst_req_1;
      type_cast_2010_inst_ack_1<= rack(0);
      type_cast_2010_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2010_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc92x_xrowx_x1_1997,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2011,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_2031_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_2031_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_2031_inst:started:   inputs: " & " type_cast_2030_wire = "& Convert_SLV_To_Hex_String(type_cast_2030_wire));
          --
        end if; 
        if type_cast_2031_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_2031_inst:finished:  outputs: " & " conv17_2032= "  & Convert_SLV_To_Hex_String(conv17_2032));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_2031_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2031_inst_req_0;
      type_cast_2031_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2031_inst_req_1;
      type_cast_2031_inst_ack_1<= rack(0);
      type_cast_2031_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2031_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2030_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2032,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_2039_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_2039_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_2039_inst:started:   inputs: " & " type_cast_2038_wire = "& Convert_SLV_To_Hex_String(type_cast_2038_wire));
          --
        end if; 
        if type_cast_2039_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_2039_inst:finished:  outputs: " & " conv104_2040= "  & Convert_SLV_To_Hex_String(conv104_2040));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_2039_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2039_inst_req_0;
      type_cast_2039_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2039_inst_req_1;
      type_cast_2039_inst_ack_1<= rack(0);
      type_cast_2039_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2039_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2038_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_2040,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator ptr_deref_1724_addr_0 flow-through 
    process(ptr_deref_1724_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1724_addr_0:flowthrough  inputs: " & " ptr_deref_1724_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1724_root_address) & "outputs: " & " ptr_deref_1724_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1724_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1724_addr_0
    process(ptr_deref_1724_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1724_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1724_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1724_base_resize flow-through 
    process(ptr_deref_1724_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1724_base_resize:flowthrough  inputs: " & " iNsTr_2_1721 = "& Convert_SLV_To_Hex_String(iNsTr_2_1721) & "outputs: " & " ptr_deref_1724_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1724_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1724_base_resize
    process(iNsTr_2_1721) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1721;
      ov := iv(6 downto 0);
      ptr_deref_1724_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1724_gather_scatter flow-through 
    process(tmp_1725) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1724_gather_scatter:flowthrough  inputs: " & " ptr_deref_1724_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1724_data_0) & "outputs: " & " tmp_1725= "  & Convert_SLV_To_Hex_String(tmp_1725));
      --
    end process; 
    -- equivalence ptr_deref_1724_gather_scatter
    process(ptr_deref_1724_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1724_data_0;
      ov(31 downto 0) := iv;
      tmp_1725 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1724_root_address_inst flow-through 
    process(ptr_deref_1724_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1724_root_address_inst:flowthrough  inputs: " & " ptr_deref_1724_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1724_resized_base_address) & "outputs: " & " ptr_deref_1724_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1724_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1724_root_address_inst
    process(ptr_deref_1724_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1724_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1724_root_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1736_addr_0 flow-through 
    process(ptr_deref_1736_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1736_addr_0:flowthrough  inputs: " & " ptr_deref_1736_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1736_root_address) & "outputs: " & " ptr_deref_1736_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1736_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1736_addr_0
    process(ptr_deref_1736_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1736_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1736_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1736_base_resize flow-through 
    process(ptr_deref_1736_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1736_base_resize:flowthrough  inputs: " & " iNsTr_3_1733 = "& Convert_SLV_To_Hex_String(iNsTr_3_1733) & "outputs: " & " ptr_deref_1736_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1736_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1736_base_resize
    process(iNsTr_3_1733) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1733;
      ov := iv(6 downto 0);
      ptr_deref_1736_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1736_gather_scatter flow-through 
    process(tmp2_1737) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1736_gather_scatter:flowthrough  inputs: " & " ptr_deref_1736_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1736_data_0) & "outputs: " & " tmp2_1737= "  & Convert_SLV_To_Hex_String(tmp2_1737));
      --
    end process; 
    -- equivalence ptr_deref_1736_gather_scatter
    process(ptr_deref_1736_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1736_data_0;
      ov(31 downto 0) := iv;
      tmp2_1737 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1736_root_address_inst flow-through 
    process(ptr_deref_1736_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1736_root_address_inst:flowthrough  inputs: " & " ptr_deref_1736_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1736_resized_base_address) & "outputs: " & " ptr_deref_1736_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1736_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1736_root_address_inst
    process(ptr_deref_1736_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1736_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1736_root_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1748_base_resize flow-through 
    process(ptr_deref_1748_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_base_resize:flowthrough  inputs: " & " iNsTr_4_1745 = "& Convert_SLV_To_Hex_String(iNsTr_4_1745) & "outputs: " & " ptr_deref_1748_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1748_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1748_base_resize
    process(iNsTr_4_1745) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1745;
      ov := iv(8 downto 0);
      ptr_deref_1748_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1748_gather_scatter flow-through 
    process(tmp5_1749) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_gather_scatter:flowthrough  inputs: " & " ptr_deref_1748_data_3 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_data_3) & " ptr_deref_1748_data_2 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_data_2) & " ptr_deref_1748_data_1 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_data_1) & " ptr_deref_1748_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_data_0) & "outputs: " & " tmp5_1749= "  & Convert_SLV_To_Hex_String(tmp5_1749));
      --
    end process; 
    -- equivalence ptr_deref_1748_gather_scatter
    process(ptr_deref_1748_data_3, ptr_deref_1748_data_2, ptr_deref_1748_data_1, ptr_deref_1748_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1748_data_3 & ptr_deref_1748_data_2 & ptr_deref_1748_data_1 & ptr_deref_1748_data_0;
      ov(31 downto 0) := iv;
      tmp5_1749 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1748_root_address_inst flow-through 
    process(ptr_deref_1748_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_root_address_inst:flowthrough  inputs: " & " ptr_deref_1748_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1748_resized_base_address) & "outputs: " & " ptr_deref_1748_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1748_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1748_root_address_inst
    process(ptr_deref_1748_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1748_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_1748_root_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1760_addr_0 flow-through 
    process(ptr_deref_1760_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1760_addr_0:flowthrough  inputs: " & " ptr_deref_1760_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1760_root_address) & "outputs: " & " ptr_deref_1760_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1760_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1760_addr_0
    process(ptr_deref_1760_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1760_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1760_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1760_base_resize flow-through 
    process(ptr_deref_1760_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1760_base_resize:flowthrough  inputs: " & " iNsTr_5_1757 = "& Convert_SLV_To_Hex_String(iNsTr_5_1757) & "outputs: " & " ptr_deref_1760_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1760_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1760_base_resize
    process(iNsTr_5_1757) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1757;
      ov := iv(6 downto 0);
      ptr_deref_1760_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1760_gather_scatter flow-through 
    process(tmp8_1761) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1760_gather_scatter:flowthrough  inputs: " & " ptr_deref_1760_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1760_data_0) & "outputs: " & " tmp8_1761= "  & Convert_SLV_To_Hex_String(tmp8_1761));
      --
    end process; 
    -- equivalence ptr_deref_1760_gather_scatter
    process(ptr_deref_1760_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1760_data_0;
      ov(31 downto 0) := iv;
      tmp8_1761 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1760_root_address_inst flow-through 
    process(ptr_deref_1760_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1760_root_address_inst:flowthrough  inputs: " & " ptr_deref_1760_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1760_resized_base_address) & "outputs: " & " ptr_deref_1760_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1760_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1760_root_address_inst
    process(ptr_deref_1760_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1760_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1760_root_address <= ov(6 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1842_branch_req_0," req0 do_while_stmt_1842_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1842_branch_ack_0," ack0 do_while_stmt_1842_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1842_branch_ack_1," ack1 do_while_stmt_1842_branch");
    do_while_stmt_1842_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2022_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1842_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1842_branch_req_0,
          ack0 => do_while_stmt_1842_branch_ack_0,
          ack1 => do_while_stmt_1842_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_2023_branch_req_0," req0 if_stmt_2023_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_2023_branch_ack_0," ack0 if_stmt_2023_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_2023_branch_ack_1," ack1 if_stmt_2023_branch");
    if_stmt_2023_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= whilex_xbody_whilex_xend_taken_2019;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2023_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2023_branch_req_0,
          ack0 => if_stmt_2023_branch_ack_0,
          ack1 => if_stmt_2023_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u16_u16_1944_inst flow-through 
    process(inc_1945) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u16_u16_1944_inst:flowthrough inputs: " & " chlx_x0_1854 = "& Convert_SLV_To_Hex_String(chlx_x0_1854) & " type_cast_1943_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1943_wire_constant) & " outputs:" & " inc_1945= "  & Convert_SLV_To_Hex_String(inc_1945));
      --
    end process; 
    -- binary operator ADD_u16_u16_1944_inst
    process(chlx_x0_1854) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chlx_x0_1854, type_cast_1943_wire_constant, tmp_var);
      inc_1945 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1965_inst flow-through 
    process(inc83x_xcolx_x1_1966) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u16_u16_1965_inst:flowthrough inputs: " & " inc83_1958 = "& Convert_SLV_To_Hex_String(inc83_1958) & " colx_x1_1949_delayed_2_0_1961 = "& Convert_SLV_To_Hex_String(colx_x1_1949_delayed_2_0_1961) & " outputs:" & " inc83x_xcolx_x1_1966= "  & Convert_SLV_To_Hex_String(inc83x_xcolx_x1_1966));
      --
    end process; 
    -- binary operator ADD_u16_u16_1965_inst
    process(inc83_1958, colx_x1_1949_delayed_2_0_1961) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc83_1958, colx_x1_1949_delayed_2_0_1961, tmp_var);
      inc83x_xcolx_x1_1966 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1996_inst flow-through 
    process(inc92x_xrowx_x1_1997) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u16_u16_1996_inst:flowthrough inputs: " & " inc92_1989 = "& Convert_SLV_To_Hex_String(inc92_1989) & " rowx_x1_1974_delayed_4_0_1992 = "& Convert_SLV_To_Hex_String(rowx_x1_1974_delayed_4_0_1992) & " outputs:" & " inc92x_xrowx_x1_1997= "  & Convert_SLV_To_Hex_String(inc92x_xrowx_x1_1997));
      --
    end process; 
    -- binary operator ADD_u16_u16_1996_inst
    process(inc92_1989, rowx_x1_1974_delayed_4_0_1992) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc92_1989, rowx_x1_1974_delayed_4_0_1992, tmp_var);
      inc92x_xrowx_x1_1997 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1816_inst flow-through 
    process(add_1817) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u32_u32_1816_inst:flowthrough inputs: " & " conv27_1794 = "& Convert_SLV_To_Hex_String(conv27_1794) & " conv14_1779 = "& Convert_SLV_To_Hex_String(conv14_1779) & " outputs:" & " add_1817= "  & Convert_SLV_To_Hex_String(add_1817));
      --
    end process; 
    -- binary operator ADD_u32_u32_1816_inst
    process(conv27_1794, conv14_1779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv27_1794, conv14_1779, tmp_var);
      add_1817 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1880_inst flow-through 
    process(add43_1881) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u32_u32_1880_inst:flowthrough inputs: " & " conv37_1867 = "& Convert_SLV_To_Hex_String(conv37_1867) & " mul42_1876 = "& Convert_SLV_To_Hex_String(mul42_1876) & " outputs:" & " add43_1881= "  & Convert_SLV_To_Hex_String(add43_1881));
      --
    end process; 
    -- binary operator ADD_u32_u32_1880_inst
    process(conv37_1867, mul42_1876) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv37_1867, mul42_1876, tmp_var);
      add43_1881 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1890_inst flow-through 
    process(add45_1891) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u32_u32_1890_inst:flowthrough inputs: " & " mul44_1886 = "& Convert_SLV_To_Hex_String(mul44_1886) & " conv33_1863 = "& Convert_SLV_To_Hex_String(conv33_1863) & " outputs:" & " add45_1891= "  & Convert_SLV_To_Hex_String(add45_1891));
      --
    end process; 
    -- binary operator ADD_u32_u32_1890_inst
    process(mul44_1886, conv33_1863) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul44_1886, conv33_1863, tmp_var);
      add45_1891 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1906_inst flow-through 
    process(add57_1907) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u32_u32_1906_inst:flowthrough inputs: " & " conv37_1867 = "& Convert_SLV_To_Hex_String(conv37_1867) & " mul56_1902 = "& Convert_SLV_To_Hex_String(mul56_1902) & " outputs:" & " add57_1907= "  & Convert_SLV_To_Hex_String(add57_1907));
      --
    end process; 
    -- binary operator ADD_u32_u32_1906_inst
    process(conv37_1867, mul56_1902) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv37_1867, mul56_1902, tmp_var);
      add57_1907 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1916_inst flow-through 
    process(add60_1917) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u32_u32_1916_inst:flowthrough inputs: " & " shl59_1912 = "& Convert_SLV_To_Hex_String(shl59_1912) & " conv33_1863 = "& Convert_SLV_To_Hex_String(conv33_1863) & " outputs:" & " add60_1917= "  & Convert_SLV_To_Hex_String(add60_1917));
      --
    end process; 
    -- binary operator ADD_u32_u32_1916_inst
    process(shl59_1912, conv33_1863) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl59_1912, conv33_1863, tmp_var);
      add60_1917 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1921_inst flow-through 
    process(add67_1922) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u32_u32_1921_inst:flowthrough inputs: " & " add60_1917 = "& Convert_SLV_To_Hex_String(add60_1917) & " conv14_1779 = "& Convert_SLV_To_Hex_String(conv14_1779) & " outputs:" & " add67_1922= "  & Convert_SLV_To_Hex_String(add67_1922));
      --
    end process; 
    -- binary operator ADD_u32_u32_1921_inst
    process(add60_1917, conv14_1779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add60_1917, conv14_1779, tmp_var);
      add67_1922 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1926_inst flow-through 
    process(add71_1927) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u32_u32_1926_inst:flowthrough inputs: " & " add60_1917 = "& Convert_SLV_To_Hex_String(add60_1917) & " conv27_1794 = "& Convert_SLV_To_Hex_String(conv27_1794) & " outputs:" & " add71_1927= "  & Convert_SLV_To_Hex_String(add71_1927));
      --
    end process; 
    -- binary operator ADD_u32_u32_1926_inst
    process(add60_1917, conv27_1794) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add60_1917, conv27_1794, tmp_var);
      add71_1927 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1931_inst flow-through 
    process(add74_1932) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ADD_u32_u32_1931_inst:flowthrough inputs: " & " add_1817 = "& Convert_SLV_To_Hex_String(add_1817) & " add60_1917 = "& Convert_SLV_To_Hex_String(add60_1917) & " outputs:" & " add74_1932= "  & Convert_SLV_To_Hex_String(add74_1932));
      --
    end process; 
    -- binary operator ADD_u32_u32_1931_inst
    process(add_1817, add60_1917) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1817, add60_1917, tmp_var);
      add74_1932 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u32_u32_1772_inst flow-through 
    process(conv12_1773) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:AND_u32_u32_1772_inst:flowthrough inputs: " & " tmp5_1749 = "& Convert_SLV_To_Hex_String(tmp5_1749) & " type_cast_1771_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1771_wire_constant) & " outputs:" & " conv12_1773= "  & Convert_SLV_To_Hex_String(conv12_1773));
      --
    end process; 
    -- binary operator AND_u32_u32_1772_inst
    process(tmp5_1749) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(tmp5_1749, type_cast_1771_wire_constant, tmp_var);
      conv12_1773 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u32_u32_1778_inst flow-through 
    process(conv14_1779) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:AND_u32_u32_1778_inst:flowthrough inputs: " & " shr_1767 = "& Convert_SLV_To_Hex_String(shr_1767) & " type_cast_1777_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1777_wire_constant) & " outputs:" & " conv14_1779= "  & Convert_SLV_To_Hex_String(conv14_1779));
      --
    end process; 
    -- binary operator AND_u32_u32_1778_inst
    process(shr_1767) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr_1767, type_cast_1777_wire_constant, tmp_var);
      conv14_1779 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u32_u32_1793_inst flow-through 
    process(conv27_1794) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:AND_u32_u32_1793_inst:flowthrough inputs: " & " mul_1784 = "& Convert_SLV_To_Hex_String(mul_1784) & " type_cast_1792_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1792_wire_constant) & " outputs:" & " conv27_1794= "  & Convert_SLV_To_Hex_String(conv27_1794));
      --
    end process; 
    -- binary operator AND_u32_u32_1793_inst
    process(mul_1784) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul_1784, type_cast_1792_wire_constant, tmp_var);
      conv27_1794 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u32_u32_1799_inst flow-through 
    process(conv39_1800) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:AND_u32_u32_1799_inst:flowthrough inputs: " & " tmp_1725 = "& Convert_SLV_To_Hex_String(tmp_1725) & " type_cast_1798_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1798_wire_constant) & " outputs:" & " conv39_1800= "  & Convert_SLV_To_Hex_String(conv39_1800));
      --
    end process; 
    -- binary operator AND_u32_u32_1799_inst
    process(tmp_1725) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(tmp_1725, type_cast_1798_wire_constant, tmp_var);
      conv39_1800 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u32_u32_1811_inst flow-through 
    process(mul58_1812) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:AND_u32_u32_1811_inst:flowthrough inputs: " & " iNsTr_8_1806 = "& Convert_SLV_To_Hex_String(iNsTr_8_1806) & " type_cast_1810_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1810_wire_constant) & " outputs:" & " mul58_1812= "  & Convert_SLV_To_Hex_String(mul58_1812));
      --
    end process; 
    -- binary operator AND_u32_u32_1811_inst
    process(iNsTr_8_1806) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_8_1806, type_cast_1810_wire_constant, tmp_var);
      mul58_1812 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u32_u32_1822_inst flow-through 
    process(conv97_1823) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:AND_u32_u32_1822_inst:flowthrough inputs: " & " tmp2_1737 = "& Convert_SLV_To_Hex_String(tmp2_1737) & " type_cast_1821_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1821_wire_constant) & " outputs:" & " conv97_1823= "  & Convert_SLV_To_Hex_String(conv97_1823));
      --
    end process; 
    -- binary operator AND_u32_u32_1822_inst
    process(tmp2_1737) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(tmp2_1737, type_cast_1821_wire_constant, tmp_var);
      conv97_1823 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u32_u1_1953_inst flow-through 
    process(cmp_1954) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:EQ_u32_u1_1953_inst:flowthrough inputs: " & " conv78_1949 = "& Convert_SLV_To_Hex_String(conv78_1949) & " conv14_1779 = "& Convert_SLV_To_Hex_String(conv14_1779) & " outputs:" & " cmp_1954= "  & Convert_SLV_To_Hex_String(cmp_1954));
      --
    end process; 
    -- binary operator EQ_u32_u1_1953_inst
    process(conv78_1949, conv14_1779) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv78_1949, conv14_1779, tmp_var);
      cmp_1954 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u32_u1_1984_inst flow-through 
    process(cmp88_1985) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:EQ_u32_u1_1984_inst:flowthrough inputs: " & " conv85_1980 = "& Convert_SLV_To_Hex_String(conv85_1980) & " conv39_1800 = "& Convert_SLV_To_Hex_String(conv39_1800) & " outputs:" & " cmp88_1985= "  & Convert_SLV_To_Hex_String(cmp88_1985));
      --
    end process; 
    -- binary operator EQ_u32_u1_1984_inst
    process(conv85_1980, conv39_1800) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv85_1980, conv39_1800, tmp_var);
      cmp88_1985 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u32_u1_2015_inst flow-through 
    process(cmp98_2016) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:EQ_u32_u1_2015_inst:flowthrough inputs: " & " conv95_2011 = "& Convert_SLV_To_Hex_String(conv95_2011) & " conv97_1823 = "& Convert_SLV_To_Hex_String(conv97_1823) & " outputs:" & " cmp98_2016= "  & Convert_SLV_To_Hex_String(cmp98_2016));
      --
    end process; 
    -- binary operator EQ_u32_u1_2015_inst
    process(conv95_2011, conv97_1823) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv95_2011, conv97_1823, tmp_var);
      cmp98_2016 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u32_u32_1766_inst flow-through 
    process(shr_1767) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:LSHR_u32_u32_1766_inst:flowthrough inputs: " & " tmp8_1761 = "& Convert_SLV_To_Hex_String(tmp8_1761) & " type_cast_1765_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1765_wire_constant) & " outputs:" & " shr_1767= "  & Convert_SLV_To_Hex_String(shr_1767));
      --
    end process; 
    -- binary operator LSHR_u32_u32_1766_inst
    process(tmp8_1761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp8_1761, type_cast_1765_wire_constant, tmp_var);
      shr_1767 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u32_u32_1805_inst flow-through 
    process(iNsTr_8_1806) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:LSHR_u32_u32_1805_inst:flowthrough inputs: " & " tmp8_1761 = "& Convert_SLV_To_Hex_String(tmp8_1761) & " type_cast_1804_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1804_wire_constant) & " outputs:" & " iNsTr_8_1806= "  & Convert_SLV_To_Hex_String(iNsTr_8_1806));
      --
    end process; 
    -- binary operator LSHR_u32_u32_1805_inst
    process(tmp8_1761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp8_1761, type_cast_1804_wire_constant, tmp_var);
      iNsTr_8_1806 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_1783_inst flow-through 
    process(mul_1784) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:MUL_u32_u32_1783_inst:flowthrough inputs: " & " conv14_1779 = "& Convert_SLV_To_Hex_String(conv14_1779) & " conv12_1773 = "& Convert_SLV_To_Hex_String(conv12_1773) & " outputs:" & " mul_1784= "  & Convert_SLV_To_Hex_String(mul_1784));
      --
    end process; 
    -- binary operator MUL_u32_u32_1783_inst
    process(conv14_1779, conv12_1773) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv14_1779, conv12_1773, tmp_var);
      mul_1784 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_1875_inst flow-through 
    process(mul42_1876) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:MUL_u32_u32_1875_inst:flowthrough inputs: " & " conv41_1871 = "& Convert_SLV_To_Hex_String(conv41_1871) & " conv39_1800 = "& Convert_SLV_To_Hex_String(conv39_1800) & " outputs:" & " mul42_1876= "  & Convert_SLV_To_Hex_String(mul42_1876));
      --
    end process; 
    -- binary operator MUL_u32_u32_1875_inst
    process(conv41_1871, conv39_1800) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv41_1871, conv39_1800, tmp_var);
      mul42_1876 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_1885_inst flow-through 
    process(mul44_1886) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:MUL_u32_u32_1885_inst:flowthrough inputs: " & " add43_1881 = "& Convert_SLV_To_Hex_String(add43_1881) & " conv14_1779 = "& Convert_SLV_To_Hex_String(conv14_1779) & " outputs:" & " mul44_1886= "  & Convert_SLV_To_Hex_String(mul44_1886));
      --
    end process; 
    -- binary operator MUL_u32_u32_1885_inst
    process(add43_1881, conv14_1779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add43_1881, conv14_1779, tmp_var);
      mul44_1886 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_1901_inst flow-through 
    process(mul56_1902) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:MUL_u32_u32_1901_inst:flowthrough inputs: " & " conv41_1871 = "& Convert_SLV_To_Hex_String(conv41_1871) & " conv12_1773 = "& Convert_SLV_To_Hex_String(conv12_1773) & " outputs:" & " mul56_1902= "  & Convert_SLV_To_Hex_String(mul56_1902));
      --
    end process; 
    -- binary operator MUL_u32_u32_1901_inst
    process(conv41_1871, conv12_1773) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv41_1871, conv12_1773, tmp_var);
      mul56_1902 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_1911_inst flow-through 
    process(shl59_1912) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:MUL_u32_u32_1911_inst:flowthrough inputs: " & " mul58_1812 = "& Convert_SLV_To_Hex_String(mul58_1812) & " add57_1907 = "& Convert_SLV_To_Hex_String(add57_1907) & " outputs:" & " shl59_1912= "  & Convert_SLV_To_Hex_String(shl59_1912));
      --
    end process; 
    -- binary operator MUL_u32_u32_1911_inst
    process(mul58_1812, add57_1907) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul58_1812, add57_1907, tmp_var);
      shl59_1912 <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_2022_inst flow-through 
    process(NOT_u1_u1_2022_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:NOT_u1_u1_2022_inst:flowthrough inputs: " & " cmp98_2016 = "& Convert_SLV_To_Hex_String(cmp98_2016) & " outputs:" & " NOT_u1_u1_2022_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_2022_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_2022_inst
    process(cmp98_2016) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp98_2016, tmp_var);
      NOT_u1_u1_2022_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator SHL_u32_u32_1896_inst flow-through 
    process(shl_1897) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:SHL_u32_u32_1896_inst:flowthrough inputs: " & " add45_1891 = "& Convert_SLV_To_Hex_String(add45_1891) & " type_cast_1895_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1895_wire_constant) & " outputs:" & " shl_1897= "  & Convert_SLV_To_Hex_String(shl_1897));
      --
    end process; 
    -- binary operator SHL_u32_u32_1896_inst
    process(add45_1891) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add45_1891, type_cast_1895_wire_constant, tmp_var);
      shl_1897 <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u64_u64_2044_inst flow-through 
    process(sub_2045) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:SUB_u64_u64_2044_inst:flowthrough inputs: " & " conv104_2040 = "& Convert_SLV_To_Hex_String(conv104_2040) & " conv17_2032 = "& Convert_SLV_To_Hex_String(conv17_2032) & " outputs:" & " sub_2045= "  & Convert_SLV_To_Hex_String(sub_2045));
      --
    end process; 
    -- binary operator SUB_u64_u64_2044_inst
    process(conv104_2040, conv17_2032) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv104_2040, conv17_2032, tmp_var);
      sub_2045 <= tmp_var; --
    end process;
    -- logger for split-operator ptr_deref_1748_addr_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1748_addr_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_addr_0:started:   inputs: " & " ptr_deref_1748_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1748_root_address) & " ptr_deref_1748_word_offset_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_word_offset_0));
          --
        end if; 
        if ptr_deref_1748_addr_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_addr_0:finished:  outputs: " & " ptr_deref_1748_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1748_word_address_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (30) : ptr_deref_1748_addr_0 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1748_root_address;
      ptr_deref_1748_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1748_addr_0_req_0;
      ptr_deref_1748_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1748_addr_0_req_1;
      ptr_deref_1748_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- logger for split-operator ptr_deref_1748_addr_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1748_addr_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_addr_1:started:   inputs: " & " ptr_deref_1748_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1748_root_address) & " ptr_deref_1748_word_offset_1 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_word_offset_1));
          --
        end if; 
        if ptr_deref_1748_addr_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_addr_1:finished:  outputs: " & " ptr_deref_1748_word_address_1= "  & Convert_SLV_To_Hex_String(ptr_deref_1748_word_address_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (31) : ptr_deref_1748_addr_1 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1748_root_address;
      ptr_deref_1748_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1748_addr_1_req_0;
      ptr_deref_1748_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1748_addr_1_req_1;
      ptr_deref_1748_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- logger for split-operator ptr_deref_1748_addr_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1748_addr_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_addr_2:started:   inputs: " & " ptr_deref_1748_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1748_root_address) & " ptr_deref_1748_word_offset_2 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_word_offset_2));
          --
        end if; 
        if ptr_deref_1748_addr_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_addr_2:finished:  outputs: " & " ptr_deref_1748_word_address_2= "  & Convert_SLV_To_Hex_String(ptr_deref_1748_word_address_2));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (32) : ptr_deref_1748_addr_2 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1748_root_address;
      ptr_deref_1748_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1748_addr_2_req_0;
      ptr_deref_1748_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1748_addr_2_req_1;
      ptr_deref_1748_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- logger for split-operator ptr_deref_1748_addr_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1748_addr_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_addr_3:started:   inputs: " & " ptr_deref_1748_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1748_root_address) & " ptr_deref_1748_word_offset_3 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_word_offset_3));
          --
        end if; 
        if ptr_deref_1748_addr_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_addr_3:finished:  outputs: " & " ptr_deref_1748_word_address_3= "  & Convert_SLV_To_Hex_String(ptr_deref_1748_word_address_3));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (33) : ptr_deref_1748_addr_3 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1748_root_address;
      ptr_deref_1748_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1748_addr_3_req_0;
      ptr_deref_1748_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1748_addr_3_req_1;
      ptr_deref_1748_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- logger for split-operator type_cast_2030_inst flow-through 
    process(type_cast_2030_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_2030_inst:flowthrough inputs: " & " call_1787 = "& Convert_SLV_To_Hex_String(call_1787) & " outputs:" & " type_cast_2030_wire= "  & Convert_SLV_To_Hex_String(type_cast_2030_wire));
      --
    end process; 
    -- unary operator type_cast_2030_inst
    process(call_1787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call_1787, tmp_var);
      type_cast_2030_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_2038_inst flow-through 
    process(type_cast_2038_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:type_cast_2038_inst:flowthrough inputs: " & " call103_2035 = "& Convert_SLV_To_Hex_String(call103_2035) & " outputs:" & " type_cast_2038_wire= "  & Convert_SLV_To_Hex_String(type_cast_2038_wire));
      --
    end process; 
    -- unary operator type_cast_2038_inst
    process(call103_2035) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call103_2035, tmp_var);
      type_cast_2038_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator ptr_deref_1724_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1724_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1724_load_0:started:   inputs: " & " ptr_deref_1724_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1724_word_address_0));
          --
        end if; 
        if ptr_deref_1724_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1724_load_0:finished:  outputs: " & " ptr_deref_1724_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1724_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_1736_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1736_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1736_load_0:started:   inputs: " & " ptr_deref_1736_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1736_word_address_0));
          --
        end if; 
        if ptr_deref_1736_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1736_load_0:finished:  outputs: " & " ptr_deref_1736_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1736_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_1760_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1760_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1760_load_0:started:   inputs: " & " ptr_deref_1760_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1760_word_address_0));
          --
        end if; 
        if ptr_deref_1760_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1760_load_0:finished:  outputs: " & " ptr_deref_1760_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1760_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : ptr_deref_1724_load_0 ptr_deref_1736_load_0 ptr_deref_1760_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1724_load_0_req_0,
        ptr_deref_1724_load_0_ack_0,
        ptr_deref_1724_load_0_req_1,
        ptr_deref_1724_load_0_ack_1,
        "ptr_deref_1724_load_0",
        "memory_space_3" ,
        ptr_deref_1724_data_0,
        ptr_deref_1724_word_address_0,
        "ptr_deref_1724_data_0",
        "ptr_deref_1724_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1736_load_0_req_0,
        ptr_deref_1736_load_0_ack_0,
        ptr_deref_1736_load_0_req_1,
        ptr_deref_1736_load_0_ack_1,
        "ptr_deref_1736_load_0",
        "memory_space_3" ,
        ptr_deref_1736_data_0,
        ptr_deref_1736_word_address_0,
        "ptr_deref_1736_data_0",
        "ptr_deref_1736_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1760_load_0_req_0,
        ptr_deref_1760_load_0_ack_0,
        ptr_deref_1760_load_0_req_1,
        ptr_deref_1760_load_0_ack_1,
        "ptr_deref_1760_load_0",
        "memory_space_3" ,
        ptr_deref_1760_data_0,
        ptr_deref_1760_word_address_0,
        "ptr_deref_1760_data_0",
        "ptr_deref_1760_word_address_0" -- 
      );
      reqL_unguarded(2) <= ptr_deref_1724_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1736_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1760_load_0_req_0;
      ptr_deref_1724_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1736_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1760_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1724_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1736_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1760_load_0_req_1;
      ptr_deref_1724_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1736_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1760_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1724_word_address_0 & ptr_deref_1736_word_address_0 & ptr_deref_1760_word_address_0;
      ptr_deref_1724_data_0 <= data_out(95 downto 64);
      ptr_deref_1736_data_0 <= data_out(63 downto 32);
      ptr_deref_1760_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator ptr_deref_1748_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1748_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_load_0:started:   inputs: " & " ptr_deref_1748_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_word_address_0));
          --
        end if; 
        if ptr_deref_1748_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_load_0:finished:  outputs: " & " ptr_deref_1748_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1748_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_1748_load_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1748_load_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_load_1:started:   inputs: " & " ptr_deref_1748_word_address_1 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_word_address_1));
          --
        end if; 
        if ptr_deref_1748_load_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_load_1:finished:  outputs: " & " ptr_deref_1748_data_1= "  & Convert_SLV_To_Hex_String(ptr_deref_1748_data_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_1748_load_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1748_load_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_load_2:started:   inputs: " & " ptr_deref_1748_word_address_2 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_word_address_2));
          --
        end if; 
        if ptr_deref_1748_load_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_load_2:finished:  outputs: " & " ptr_deref_1748_data_2= "  & Convert_SLV_To_Hex_String(ptr_deref_1748_data_2));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_1748_load_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1748_load_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_load_3:started:   inputs: " & " ptr_deref_1748_word_address_3 = "& Convert_SLV_To_Hex_String(ptr_deref_1748_word_address_3));
          --
        end if; 
        if ptr_deref_1748_load_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:ptr_deref_1748_load_3:finished:  outputs: " & " ptr_deref_1748_data_3= "  & Convert_SLV_To_Hex_String(ptr_deref_1748_data_3));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (1) : ptr_deref_1748_load_0 ptr_deref_1748_load_1 ptr_deref_1748_load_2 ptr_deref_1748_load_3 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1748_load_0_req_0,
        ptr_deref_1748_load_0_ack_0,
        ptr_deref_1748_load_0_req_1,
        ptr_deref_1748_load_0_ack_1,
        "ptr_deref_1748_load_0",
        "memory_space_4" ,
        ptr_deref_1748_data_0,
        ptr_deref_1748_word_address_0,
        "ptr_deref_1748_data_0",
        "ptr_deref_1748_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1748_load_1_req_0,
        ptr_deref_1748_load_1_ack_0,
        ptr_deref_1748_load_1_req_1,
        ptr_deref_1748_load_1_ack_1,
        "ptr_deref_1748_load_1",
        "memory_space_4" ,
        ptr_deref_1748_data_1,
        ptr_deref_1748_word_address_1,
        "ptr_deref_1748_data_1",
        "ptr_deref_1748_word_address_1" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1748_load_2_req_0,
        ptr_deref_1748_load_2_ack_0,
        ptr_deref_1748_load_2_req_1,
        ptr_deref_1748_load_2_ack_1,
        "ptr_deref_1748_load_2",
        "memory_space_4" ,
        ptr_deref_1748_data_2,
        ptr_deref_1748_word_address_2,
        "ptr_deref_1748_data_2",
        "ptr_deref_1748_word_address_2" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1748_load_3_req_0,
        ptr_deref_1748_load_3_ack_0,
        ptr_deref_1748_load_3_req_1,
        ptr_deref_1748_load_3_ack_1,
        "ptr_deref_1748_load_3",
        "memory_space_4" ,
        ptr_deref_1748_data_3,
        ptr_deref_1748_word_address_3,
        "ptr_deref_1748_data_3",
        "ptr_deref_1748_word_address_3" -- 
      );
      reqL_unguarded(3) <= ptr_deref_1748_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1748_load_1_req_0;
      reqL_unguarded(1) <= ptr_deref_1748_load_2_req_0;
      reqL_unguarded(0) <= ptr_deref_1748_load_3_req_0;
      ptr_deref_1748_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1748_load_1_ack_0 <= ackL_unguarded(2);
      ptr_deref_1748_load_2_ack_0 <= ackL_unguarded(1);
      ptr_deref_1748_load_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_1748_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1748_load_1_req_1;
      reqR_unguarded(1) <= ptr_deref_1748_load_2_req_1;
      reqR_unguarded(0) <= ptr_deref_1748_load_3_req_1;
      ptr_deref_1748_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1748_load_1_ack_1 <= ackR_unguarded(2);
      ptr_deref_1748_load_2_ack_1 <= ackR_unguarded(1);
      ptr_deref_1748_load_3_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1748_word_address_0 & ptr_deref_1748_word_address_1 & ptr_deref_1748_word_address_2 & ptr_deref_1748_word_address_3;
      ptr_deref_1748_data_0 <= data_out(31 downto 24);
      ptr_deref_1748_data_1 <= data_out(23 downto 16);
      ptr_deref_1748_data_2 <= data_out(15 downto 8);
      ptr_deref_1748_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 9,
        num_reqs => 4,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(8 downto 0),
          mtag => memory_space_4_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 8,
        num_reqs => 4,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(7 downto 0),
          mtag => memory_space_4_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- logger for split-operator WPIPE_elapsed_time_pipe_2046_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_elapsed_time_pipe_2046_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:WPIPE_elapsed_time_pipe_2046_inst:started:   PipeWrite to elapsed_time_pipe inputs: " & " sub_2045 = "& Convert_SLV_To_Hex_String(sub_2045));
          --
        end if; 
        if WPIPE_elapsed_time_pipe_2046_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:WPIPE_elapsed_time_pipe_2046_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_2046_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_2046_inst_req_0;
      WPIPE_elapsed_time_pipe_2046_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_2046_inst_req_1;
      WPIPE_elapsed_time_pipe_2046_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_2045;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_1712_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1712_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:call_stmt_1712_call:started:  Call to module testConfigure inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if call_stmt_1712_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:call_stmt_1712_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1712_call 
    testConfigure_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1712_call_req_0;
      call_stmt_1712_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1712_call_req_1;
      call_stmt_1712_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_1787_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1787_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:call_stmt_1787_call:started:  Call to module timer inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if call_stmt_1787_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:call_stmt_1787_call:finished:  outputs: " & " call_1787= "  & Convert_SLV_To_Hex_String(call_1787));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_2035_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_2035_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:call_stmt_2035_call:started:  Call to module timer inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if call_stmt_2035_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:call_stmt_2035_call:finished:  outputs: " & " call103_2035= "  & Convert_SLV_To_Hex_String(call103_2035));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_1787_call call_stmt_2035_call 
    timer_call_group_1: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1787_call_req_0;
      reqL_unguarded(0) <= call_stmt_2035_call_req_0;
      call_stmt_1787_call_ack_0 <= ackL_unguarded(1);
      call_stmt_2035_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1787_call_req_1;
      reqR_unguarded(0) <= call_stmt_2035_call_req_1;
      call_stmt_1787_call_ack_1 <= ackR_unguarded(1);
      call_stmt_2035_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_1_gI: SplitGuardInterface generic map(name => "timer_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_1787 <= data_out(127 downto 64);
      call103_2035 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_1939_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1939_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:call_stmt_1939_call:started:  Call to module maxPool4 inputs: " & " shl_1897 = "& Convert_SLV_To_Hex_String(shl_1897) & " add60_1917 = "& Convert_SLV_To_Hex_String(add60_1917) & " add67_1922 = "& Convert_SLV_To_Hex_String(add67_1922) & " add71_1927 = "& Convert_SLV_To_Hex_String(add71_1927) & " add74_1932 = "& Convert_SLV_To_Hex_String(add74_1932));
          --
        end if; 
        if call_stmt_1939_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:call_stmt_1939_call:finished:  outputs: " & " call75_1939= "  & Convert_SLV_To_Hex_String(call75_1939));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_1939_call 
    maxPool4_call_group_2: Block -- 
      signal data_in: std_logic_vector(159 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 17);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1939_call_req_0;
      call_stmt_1939_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1939_call_req_1;
      call_stmt_1939_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      maxPool4_call_group_2_gI: SplitGuardInterface generic map(name => "maxPool4_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= shl_1897 & add60_1917 & add67_1922 & add71_1927 & add74_1932;
      call75_1939 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 160,
        owidth => 160,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => maxPool4_call_reqs(0),
          ackR => maxPool4_call_acks(0),
          dataR => maxPool4_call_data(159 downto 0),
          tagR => maxPool4_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => maxPool4_return_acks(0), -- cross-over
          ackL => maxPool4_return_reqs(0), -- cross-over
          dataL => maxPool4_return_data(7 downto 0),
          tagL => maxPool4_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- logger for split-operator call_stmt_2050_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_2050_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:call_stmt_2050_call:started:  Call to module sendB inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if call_stmt_2050_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool3D:DP:call_stmt_2050_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (3) : call_stmt_2050_call 
    sendB_call_group_3: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2050_call_req_0;
      call_stmt_2050_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2050_call_req_1;
      call_stmt_2050_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendB_call_group_3_gI: SplitGuardInterface generic map(name => "sendB_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendB_call_reqs(0),
          ackR => sendB_call_acks(0),
          tagR => sendB_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendB_return_acks(0), -- cross-over
          ackL => sendB_return_reqs(0), -- cross-over
          tagL => sendB_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end maxPool3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool4 is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(31 downto 0);
    addr1 : in  std_logic_vector(31 downto 0);
    addr2 : in  std_logic_vector(31 downto 0);
    addr3 : in  std_logic_vector(31 downto 0);
    addr4 : in  std_logic_vector(31 downto 0);
    output : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool4;
architecture maxPool4_arch of maxPool4 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 160)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(31 downto 0);
  signal addr_update_enable: Boolean;
  signal addr1_buffer :  std_logic_vector(31 downto 0);
  signal addr1_update_enable: Boolean;
  signal addr2_buffer :  std_logic_vector(31 downto 0);
  signal addr2_update_enable: Boolean;
  signal addr3_buffer :  std_logic_vector(31 downto 0);
  signal addr3_update_enable: Boolean;
  signal addr4_buffer :  std_logic_vector(31 downto 0);
  signal addr4_update_enable: Boolean;
  -- output port buffer signals
  signal output_buffer :  std_logic_vector(7 downto 0);
  signal output_update_enable: Boolean;
  signal maxPool4_CP_1841_start: Boolean;
  signal maxPool4_CP_1841_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal slice_617_inst_ack_0 : boolean;
  signal array_obj_ref_422_index_offset_req_1 : boolean;
  signal slice_581_inst_req_1 : boolean;
  signal slice_589_inst_ack_0 : boolean;
  signal array_obj_ref_422_index_offset_req_0 : boolean;
  signal slice_581_inst_req_0 : boolean;
  signal slice_545_inst_ack_0 : boolean;
  signal slice_589_inst_req_0 : boolean;
  signal array_obj_ref_415_index_offset_req_0 : boolean;
  signal array_obj_ref_415_index_offset_ack_0 : boolean;
  signal slice_545_inst_req_0 : boolean;
  signal addr_of_423_final_reg_req_0 : boolean;
  signal array_obj_ref_422_index_offset_ack_1 : boolean;
  signal slice_581_inst_ack_0 : boolean;
  signal slice_541_inst_req_1 : boolean;
  signal slice_581_inst_ack_1 : boolean;
  signal addr_of_423_final_reg_ack_1 : boolean;
  signal slice_585_inst_ack_0 : boolean;
  signal slice_541_inst_req_0 : boolean;
  signal addr_of_416_final_reg_ack_1 : boolean;
  signal array_obj_ref_422_index_offset_ack_0 : boolean;
  signal array_obj_ref_415_index_offset_ack_1 : boolean;
  signal slice_605_inst_ack_0 : boolean;
  signal array_obj_ref_415_index_offset_req_1 : boolean;
  signal slice_621_inst_req_1 : boolean;
  signal slice_585_inst_req_0 : boolean;
  signal addr_of_423_final_reg_ack_0 : boolean;
  signal slice_553_inst_req_0 : boolean;
  signal array_obj_ref_429_index_offset_req_0 : boolean;
  signal slice_617_inst_req_0 : boolean;
  signal slice_561_inst_req_1 : boolean;
  signal array_obj_ref_429_index_offset_ack_0 : boolean;
  signal addr_of_423_final_reg_req_1 : boolean;
  signal array_obj_ref_429_index_offset_req_1 : boolean;
  signal slice_577_inst_req_1 : boolean;
  signal array_obj_ref_429_index_offset_ack_1 : boolean;
  signal slice_597_inst_ack_0 : boolean;
  signal slice_541_inst_ack_1 : boolean;
  signal addr_of_416_final_reg_req_0 : boolean;
  signal array_obj_ref_436_index_offset_req_1 : boolean;
  signal array_obj_ref_436_index_offset_ack_1 : boolean;
  signal slice_585_inst_ack_1 : boolean;
  signal array_obj_ref_436_index_offset_req_0 : boolean;
  signal slice_549_inst_ack_1 : boolean;
  signal slice_565_inst_req_1 : boolean;
  signal slice_561_inst_ack_0 : boolean;
  signal slice_549_inst_req_1 : boolean;
  signal addr_of_416_final_reg_ack_0 : boolean;
  signal slice_597_inst_req_0 : boolean;
  signal slice_541_inst_ack_0 : boolean;
  signal slice_605_inst_req_0 : boolean;
  signal array_obj_ref_436_index_offset_ack_0 : boolean;
  signal slice_553_inst_ack_1 : boolean;
  signal addr_of_416_final_reg_req_1 : boolean;
  signal slice_605_inst_req_1 : boolean;
  signal slice_601_inst_req_1 : boolean;
  signal slice_613_inst_ack_0 : boolean;
  signal ptr_deref_441_load_0_req_0 : boolean;
  signal slice_577_inst_ack_0 : boolean;
  signal ptr_deref_441_load_0_ack_0 : boolean;
  signal slice_537_inst_ack_1 : boolean;
  signal slice_593_inst_ack_1 : boolean;
  signal slice_613_inst_ack_1 : boolean;
  signal slice_593_inst_req_1 : boolean;
  signal slice_553_inst_req_1 : boolean;
  signal slice_593_inst_req_0 : boolean;
  signal ptr_deref_441_load_0_ack_1 : boolean;
  signal slice_601_inst_ack_1 : boolean;
  signal slice_577_inst_req_0 : boolean;
  signal slice_613_inst_req_0 : boolean;
  signal slice_577_inst_ack_1 : boolean;
  signal addr_of_430_final_reg_ack_1 : boolean;
  signal addr_of_437_final_reg_ack_1 : boolean;
  signal slice_561_inst_req_0 : boolean;
  signal addr_of_430_final_reg_req_1 : boolean;
  signal slice_605_inst_ack_1 : boolean;
  signal slice_593_inst_ack_0 : boolean;
  signal addr_of_430_final_reg_ack_0 : boolean;
  signal ptr_deref_441_load_0_req_1 : boolean;
  signal slice_621_inst_req_0 : boolean;
  signal slice_585_inst_req_1 : boolean;
  signal addr_of_430_final_reg_req_0 : boolean;
  signal addr_of_437_final_reg_req_0 : boolean;
  signal addr_of_437_final_reg_ack_0 : boolean;
  signal slice_609_inst_ack_1 : boolean;
  signal slice_609_inst_req_1 : boolean;
  signal addr_of_437_final_reg_req_1 : boolean;
  signal slice_553_inst_ack_0 : boolean;
  signal slice_601_inst_ack_0 : boolean;
  signal slice_601_inst_req_0 : boolean;
  signal slice_621_inst_ack_1 : boolean;
  signal slice_613_inst_req_1 : boolean;
  signal slice_621_inst_ack_0 : boolean;
  signal slice_609_inst_ack_0 : boolean;
  signal slice_537_inst_req_1 : boolean;
  signal slice_557_inst_ack_1 : boolean;
  signal ptr_deref_445_load_0_req_0 : boolean;
  signal ptr_deref_445_load_0_ack_0 : boolean;
  signal slice_557_inst_req_1 : boolean;
  signal ptr_deref_445_load_0_req_1 : boolean;
  signal ptr_deref_445_load_0_ack_1 : boolean;
  signal slice_609_inst_req_0 : boolean;
  signal slice_573_inst_ack_1 : boolean;
  signal slice_573_inst_req_1 : boolean;
  signal slice_549_inst_ack_0 : boolean;
  signal slice_549_inst_req_0 : boolean;
  signal slice_573_inst_ack_0 : boolean;
  signal slice_573_inst_req_0 : boolean;
  signal slice_569_inst_ack_1 : boolean;
  signal slice_569_inst_req_1 : boolean;
  signal slice_617_inst_ack_1 : boolean;
  signal slice_537_inst_ack_0 : boolean;
  signal ptr_deref_449_load_0_req_0 : boolean;
  signal ptr_deref_449_load_0_ack_0 : boolean;
  signal slice_537_inst_req_0 : boolean;
  signal slice_557_inst_ack_0 : boolean;
  signal ptr_deref_449_load_0_req_1 : boolean;
  signal slice_569_inst_ack_0 : boolean;
  signal ptr_deref_449_load_0_ack_1 : boolean;
  signal slice_569_inst_req_0 : boolean;
  signal slice_617_inst_req_1 : boolean;
  signal slice_565_inst_ack_1 : boolean;
  signal slice_625_inst_req_0 : boolean;
  signal slice_589_inst_ack_1 : boolean;
  signal slice_565_inst_ack_0 : boolean;
  signal slice_565_inst_req_0 : boolean;
  signal slice_589_inst_req_1 : boolean;
  signal slice_557_inst_req_0 : boolean;
  signal ptr_deref_453_load_0_req_0 : boolean;
  signal ptr_deref_453_load_0_ack_0 : boolean;
  signal ptr_deref_453_load_0_req_1 : boolean;
  signal ptr_deref_453_load_0_ack_1 : boolean;
  signal slice_545_inst_ack_1 : boolean;
  signal slice_597_inst_ack_1 : boolean;
  signal slice_545_inst_req_1 : boolean;
  signal slice_561_inst_ack_1 : boolean;
  signal slice_597_inst_req_1 : boolean;
  signal slice_457_inst_req_0 : boolean;
  signal slice_457_inst_ack_0 : boolean;
  signal slice_457_inst_req_1 : boolean;
  signal slice_457_inst_ack_1 : boolean;
  signal W_myptr6_1382_delayed_8_0_1385_inst_req_1 : boolean;
  signal slice_461_inst_req_0 : boolean;
  signal slice_461_inst_ack_0 : boolean;
  signal array_obj_ref_1408_index_offset_ack_1 : boolean;
  signal slice_461_inst_req_1 : boolean;
  signal slice_461_inst_ack_1 : boolean;
  signal W_myptr6_1382_delayed_8_0_1385_inst_ack_1 : boolean;
  signal slice_465_inst_req_0 : boolean;
  signal slice_465_inst_ack_0 : boolean;
  signal slice_465_inst_req_1 : boolean;
  signal slice_465_inst_ack_1 : boolean;
  signal slice_469_inst_req_0 : boolean;
  signal slice_469_inst_ack_0 : boolean;
  signal slice_469_inst_req_1 : boolean;
  signal slice_469_inst_ack_1 : boolean;
  signal slice_473_inst_req_0 : boolean;
  signal slice_473_inst_ack_0 : boolean;
  signal slice_473_inst_req_1 : boolean;
  signal slice_473_inst_ack_1 : boolean;
  signal slice_477_inst_req_0 : boolean;
  signal slice_477_inst_ack_0 : boolean;
  signal slice_477_inst_req_1 : boolean;
  signal slice_477_inst_ack_1 : boolean;
  signal slice_481_inst_req_0 : boolean;
  signal slice_481_inst_ack_0 : boolean;
  signal slice_481_inst_req_1 : boolean;
  signal slice_481_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1400_inst_req_0 : boolean;
  signal array_obj_ref_1408_index_offset_req_1 : boolean;
  signal CONCAT_u32_u64_1400_inst_ack_0 : boolean;
  signal slice_485_inst_req_0 : boolean;
  signal slice_485_inst_ack_0 : boolean;
  signal slice_485_inst_req_1 : boolean;
  signal slice_485_inst_ack_1 : boolean;
  signal slice_489_inst_req_0 : boolean;
  signal slice_489_inst_ack_0 : boolean;
  signal slice_489_inst_req_1 : boolean;
  signal slice_489_inst_ack_1 : boolean;
  signal slice_493_inst_req_0 : boolean;
  signal slice_493_inst_ack_0 : boolean;
  signal slice_493_inst_req_1 : boolean;
  signal slice_493_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1400_inst_req_1 : boolean;
  signal W_myptr7_1405_delayed_8_0_1411_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1400_inst_ack_1 : boolean;
  signal slice_497_inst_req_0 : boolean;
  signal slice_497_inst_ack_0 : boolean;
  signal slice_497_inst_req_1 : boolean;
  signal slice_497_inst_ack_1 : boolean;
  signal slice_501_inst_req_0 : boolean;
  signal slice_501_inst_ack_0 : boolean;
  signal slice_501_inst_req_1 : boolean;
  signal slice_501_inst_ack_1 : boolean;
  signal slice_505_inst_req_0 : boolean;
  signal slice_505_inst_ack_0 : boolean;
  signal slice_505_inst_req_1 : boolean;
  signal slice_505_inst_ack_1 : boolean;
  signal slice_509_inst_req_0 : boolean;
  signal slice_509_inst_ack_0 : boolean;
  signal slice_509_inst_req_1 : boolean;
  signal slice_509_inst_ack_1 : boolean;
  signal slice_513_inst_req_0 : boolean;
  signal slice_513_inst_ack_0 : boolean;
  signal slice_513_inst_req_1 : boolean;
  signal slice_513_inst_ack_1 : boolean;
  signal slice_517_inst_req_0 : boolean;
  signal slice_517_inst_ack_0 : boolean;
  signal slice_517_inst_req_1 : boolean;
  signal slice_517_inst_ack_1 : boolean;
  signal slice_521_inst_req_0 : boolean;
  signal slice_521_inst_ack_0 : boolean;
  signal slice_521_inst_req_1 : boolean;
  signal slice_521_inst_ack_1 : boolean;
  signal slice_525_inst_req_0 : boolean;
  signal slice_525_inst_ack_0 : boolean;
  signal slice_525_inst_req_1 : boolean;
  signal slice_525_inst_ack_1 : boolean;
  signal slice_529_inst_req_0 : boolean;
  signal slice_529_inst_ack_0 : boolean;
  signal slice_529_inst_req_1 : boolean;
  signal slice_529_inst_ack_1 : boolean;
  signal slice_533_inst_req_0 : boolean;
  signal slice_533_inst_ack_0 : boolean;
  signal slice_533_inst_req_1 : boolean;
  signal slice_533_inst_ack_1 : boolean;
  signal slice_705_inst_req_1 : boolean;
  signal slice_705_inst_ack_1 : boolean;
  signal slice_625_inst_ack_0 : boolean;
  signal slice_625_inst_req_1 : boolean;
  signal slice_625_inst_ack_1 : boolean;
  signal W_myptr6_1382_delayed_8_0_1385_inst_ack_0 : boolean;
  signal addr_of_1409_final_reg_ack_1 : boolean;
  signal W_myptr6_1382_delayed_8_0_1385_inst_req_0 : boolean;
  signal slice_629_inst_req_0 : boolean;
  signal slice_629_inst_ack_0 : boolean;
  signal slice_629_inst_req_1 : boolean;
  signal slice_629_inst_ack_1 : boolean;
  signal addr_of_1409_final_reg_req_1 : boolean;
  signal ptr_deref_1363_store_0_ack_1 : boolean;
  signal CONCAT_u32_u64_1426_inst_ack_1 : boolean;
  signal slice_633_inst_req_0 : boolean;
  signal slice_633_inst_ack_0 : boolean;
  signal ptr_deref_1363_store_0_req_1 : boolean;
  signal CONCAT_u32_u64_1426_inst_req_1 : boolean;
  signal slice_633_inst_req_1 : boolean;
  signal slice_633_inst_ack_1 : boolean;
  signal array_obj_ref_1408_index_offset_ack_0 : boolean;
  signal ptr_deref_1389_store_0_ack_1 : boolean;
  signal slice_637_inst_req_0 : boolean;
  signal ptr_deref_1389_store_0_req_1 : boolean;
  signal slice_637_inst_ack_0 : boolean;
  signal slice_637_inst_req_1 : boolean;
  signal slice_637_inst_ack_1 : boolean;
  signal addr_of_1383_final_reg_ack_1 : boolean;
  signal array_obj_ref_1408_index_offset_req_0 : boolean;
  signal addr_of_1383_final_reg_req_1 : boolean;
  signal CONCAT_u32_u64_1426_inst_ack_0 : boolean;
  signal slice_641_inst_req_0 : boolean;
  signal slice_641_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1426_inst_req_0 : boolean;
  signal slice_641_inst_req_1 : boolean;
  signal slice_641_inst_ack_1 : boolean;
  signal addr_of_1383_final_reg_ack_0 : boolean;
  signal addr_of_1383_final_reg_req_0 : boolean;
  signal slice_645_inst_req_0 : boolean;
  signal slice_645_inst_ack_0 : boolean;
  signal ptr_deref_1363_store_0_ack_0 : boolean;
  signal slice_645_inst_req_1 : boolean;
  signal slice_645_inst_ack_1 : boolean;
  signal ptr_deref_1363_store_0_req_0 : boolean;
  signal addr_of_1409_final_reg_ack_0 : boolean;
  signal ptr_deref_1389_store_0_ack_0 : boolean;
  signal slice_649_inst_req_0 : boolean;
  signal ptr_deref_1389_store_0_req_0 : boolean;
  signal slice_649_inst_ack_0 : boolean;
  signal slice_649_inst_req_1 : boolean;
  signal slice_649_inst_ack_1 : boolean;
  signal addr_of_1409_final_reg_req_0 : boolean;
  signal slice_653_inst_req_0 : boolean;
  signal slice_653_inst_ack_0 : boolean;
  signal slice_653_inst_req_1 : boolean;
  signal slice_653_inst_ack_1 : boolean;
  signal array_obj_ref_1382_index_offset_ack_1 : boolean;
  signal array_obj_ref_1382_index_offset_req_1 : boolean;
  signal W_myptr7_1405_delayed_8_0_1411_inst_ack_1 : boolean;
  signal slice_657_inst_req_0 : boolean;
  signal slice_657_inst_ack_0 : boolean;
  signal W_myptr7_1405_delayed_8_0_1411_inst_req_1 : boolean;
  signal slice_657_inst_req_1 : boolean;
  signal slice_657_inst_ack_1 : boolean;
  signal array_obj_ref_1382_index_offset_ack_0 : boolean;
  signal slice_661_inst_req_0 : boolean;
  signal slice_661_inst_ack_0 : boolean;
  signal slice_661_inst_req_1 : boolean;
  signal slice_661_inst_ack_1 : boolean;
  signal array_obj_ref_1382_index_offset_req_0 : boolean;
  signal W_myptr7_1405_delayed_8_0_1411_inst_ack_0 : boolean;
  signal slice_665_inst_req_0 : boolean;
  signal slice_665_inst_ack_0 : boolean;
  signal slice_665_inst_req_1 : boolean;
  signal slice_665_inst_ack_1 : boolean;
  signal slice_669_inst_req_0 : boolean;
  signal slice_669_inst_ack_0 : boolean;
  signal slice_669_inst_req_1 : boolean;
  signal slice_669_inst_ack_1 : boolean;
  signal slice_673_inst_req_0 : boolean;
  signal slice_673_inst_ack_0 : boolean;
  signal slice_673_inst_req_1 : boolean;
  signal slice_673_inst_ack_1 : boolean;
  signal slice_677_inst_req_0 : boolean;
  signal slice_677_inst_ack_0 : boolean;
  signal slice_677_inst_req_1 : boolean;
  signal slice_677_inst_ack_1 : boolean;
  signal slice_681_inst_req_0 : boolean;
  signal slice_681_inst_ack_0 : boolean;
  signal slice_681_inst_req_1 : boolean;
  signal slice_681_inst_ack_1 : boolean;
  signal slice_685_inst_req_0 : boolean;
  signal slice_685_inst_ack_0 : boolean;
  signal slice_685_inst_req_1 : boolean;
  signal slice_685_inst_ack_1 : boolean;
  signal slice_689_inst_req_0 : boolean;
  signal slice_689_inst_ack_0 : boolean;
  signal slice_689_inst_req_1 : boolean;
  signal slice_689_inst_ack_1 : boolean;
  signal slice_693_inst_req_0 : boolean;
  signal slice_693_inst_ack_0 : boolean;
  signal slice_693_inst_req_1 : boolean;
  signal slice_693_inst_ack_1 : boolean;
  signal slice_697_inst_req_0 : boolean;
  signal slice_697_inst_ack_0 : boolean;
  signal slice_697_inst_req_1 : boolean;
  signal slice_697_inst_ack_1 : boolean;
  signal slice_701_inst_req_0 : boolean;
  signal slice_701_inst_ack_0 : boolean;
  signal slice_701_inst_req_1 : boolean;
  signal slice_701_inst_ack_1 : boolean;
  signal slice_705_inst_req_0 : boolean;
  signal slice_705_inst_ack_0 : boolean;
  signal slice_709_inst_req_0 : boolean;
  signal slice_709_inst_ack_0 : boolean;
  signal slice_709_inst_req_1 : boolean;
  signal slice_709_inst_ack_1 : boolean;
  signal array_obj_ref_1356_index_offset_req_0 : boolean;
  signal array_obj_ref_1356_index_offset_ack_0 : boolean;
  signal array_obj_ref_1356_index_offset_req_1 : boolean;
  signal array_obj_ref_1356_index_offset_ack_1 : boolean;
  signal addr_of_1357_final_reg_req_0 : boolean;
  signal addr_of_1357_final_reg_ack_0 : boolean;
  signal addr_of_1357_final_reg_req_1 : boolean;
  signal addr_of_1357_final_reg_ack_1 : boolean;
  signal W_myptr5_1359_delayed_8_0_1359_inst_req_0 : boolean;
  signal W_myptr5_1359_delayed_8_0_1359_inst_ack_0 : boolean;
  signal W_myptr5_1359_delayed_8_0_1359_inst_req_1 : boolean;
  signal W_myptr5_1359_delayed_8_0_1359_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1374_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1374_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1374_inst_req_1 : boolean;
  signal CONCAT_u32_u64_1374_inst_ack_1 : boolean;
  signal ptr_deref_1415_store_0_req_0 : boolean;
  signal ptr_deref_1415_store_0_ack_0 : boolean;
  signal ptr_deref_1415_store_0_req_1 : boolean;
  signal ptr_deref_1415_store_0_ack_1 : boolean;
  signal array_obj_ref_1434_index_offset_req_0 : boolean;
  signal array_obj_ref_1434_index_offset_ack_0 : boolean;
  signal array_obj_ref_1434_index_offset_req_1 : boolean;
  signal array_obj_ref_1434_index_offset_ack_1 : boolean;
  signal addr_of_1435_final_reg_req_0 : boolean;
  signal addr_of_1435_final_reg_ack_0 : boolean;
  signal addr_of_1435_final_reg_req_1 : boolean;
  signal addr_of_1435_final_reg_ack_1 : boolean;
  signal W_myptr8_1428_delayed_8_0_1437_inst_req_0 : boolean;
  signal W_myptr8_1428_delayed_8_0_1437_inst_ack_0 : boolean;
  signal W_myptr8_1428_delayed_8_0_1437_inst_req_1 : boolean;
  signal W_myptr8_1428_delayed_8_0_1437_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1452_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1452_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1452_inst_req_1 : boolean;
  signal CONCAT_u32_u64_1452_inst_ack_1 : boolean;
  signal ptr_deref_1441_store_0_req_0 : boolean;
  signal ptr_deref_1441_store_0_ack_0 : boolean;
  signal ptr_deref_1441_store_0_req_1 : boolean;
  signal ptr_deref_1441_store_0_ack_1 : boolean;
  signal type_cast_1456_inst_req_0 : boolean;
  signal type_cast_1456_inst_ack_0 : boolean;
  signal type_cast_1456_inst_req_1 : boolean;
  signal type_cast_1456_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool4_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 160) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= addr1;
  addr1_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(95 downto 64) <= addr2;
  addr2_buffer <= in_buffer_data_out(95 downto 64);
  in_buffer_data_in(127 downto 96) <= addr3;
  addr3_buffer <= in_buffer_data_out(127 downto 96);
  in_buffer_data_in(159 downto 128) <= addr4;
  addr4_buffer <= in_buffer_data_out(159 downto 128);
  in_buffer_data_in(tag_length + 159 downto 160) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 159 downto 160);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1,6 => 15);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 15);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= addr_update_enable & addr1_update_enable & addr2_update_enable & addr3_update_enable & addr4_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool4_CP_1841_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool4_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= output_buffer;
  output <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_1841_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  output_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "output_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_output_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => output_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool4_CP_1841_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_1841_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,maxPool4_CP_1841_start,"maxPool4 cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,maxPool4_CP_1841_symbol, "maxPool4 cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool4_CP_1841: Block -- control-path 
    signal maxPool4_CP_1841_elements: BooleanArray(398 downto 0);
    -- 
  begin -- 
    maxPool4_CP_1841_elements(0) <= maxPool4_CP_1841_start;
    maxPool4_CP_1841_symbol <= maxPool4_CP_1841_elements(398);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	11 
    -- CP-element group 1: 	16 
    -- CP-element group 1: 	17 
    -- CP-element group 1: 	18 
    -- CP-element group 1: 	23 
    -- CP-element group 1: 	24 
    -- CP-element group 1: 	25 
    -- CP-element group 1: 	30 
    -- CP-element group 1: 	31 
    -- CP-element group 1: 	32 
    -- CP-element group 1: 	309 
    -- CP-element group 1: 	310 
    -- CP-element group 1: 	311 
    -- CP-element group 1: 	328 
    -- CP-element group 1: 	329 
    -- CP-element group 1: 	330 
    -- CP-element group 1: 	347 
    -- CP-element group 1: 	348 
    -- CP-element group 1: 	349 
    -- CP-element group 1: 	366 
    -- CP-element group 1: 	367 
    -- CP-element group 1: 	368 
    -- CP-element group 1:  members (105) 
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_resized_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_computed_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_computed_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_computed_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_resized_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_resized_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_computed_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_index_resized_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_resized_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_computed_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_computed_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_resized_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_resized_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_computed_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_resized_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_computed_1
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_final_index_sum_regn_Sample/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_415_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_422_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_429_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_436_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1356_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1382_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1408_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1434_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(1), ack => array_obj_ref_415_index_offset_req_0); -- 
    req_1929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(1), ack => array_obj_ref_422_index_offset_req_0); -- 
    req_1975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(1), ack => array_obj_ref_429_index_offset_req_0); -- 
    req_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(1), ack => array_obj_ref_436_index_offset_req_0); -- 
    req_3163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(1), ack => array_obj_ref_1356_index_offset_req_0); -- 
    req_3287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(1), ack => array_obj_ref_1382_index_offset_req_0); -- 
    req_3411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(1), ack => array_obj_ref_1408_index_offset_req_0); -- 
    req_3535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(1), ack => array_obj_ref_1434_index_offset_req_0); -- 
    maxPool4_CP_1841_elements(1) <= maxPool4_CP_1841_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	311 
    -- CP-element group 2: 	330 
    -- CP-element group 2: 	349 
    -- CP-element group 2: 	368 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	392 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_417_to_assign_stmt_1457/addr_update_enable_out
      -- CP-element group 2: 	 assign_stmt_417_to_assign_stmt_1457/addr_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(311) & maxPool4_CP_1841_elements(330) & maxPool4_CP_1841_elements(349) & maxPool4_CP_1841_elements(368);
      gj_maxPool4_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	11 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	393 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_417_to_assign_stmt_1457/addr1_update_enable_out
      -- CP-element group 3: 	 assign_stmt_417_to_assign_stmt_1457/addr1_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_1841_elements(11);
      gj_maxPool4_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	18 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	394 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_417_to_assign_stmt_1457/addr2_update_enable_out
      -- CP-element group 4: 	 assign_stmt_417_to_assign_stmt_1457/addr2_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_1841_elements(18);
      gj_maxPool4_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	25 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	395 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_417_to_assign_stmt_1457/addr3_update_enable_out
      -- CP-element group 5: 	 assign_stmt_417_to_assign_stmt_1457/addr3_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_1841_elements(25);
      gj_maxPool4_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	32 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	396 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_417_to_assign_stmt_1457/addr4_update_enable_out
      -- CP-element group 6: 	 assign_stmt_417_to_assign_stmt_1457/addr4_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_1841_elements(32);
      gj_maxPool4_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	397 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	385 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_417_to_assign_stmt_1457/output_update_enable_in
      -- CP-element group 7: 	 assign_stmt_417_to_assign_stmt_1457/output_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_CP_1841_elements(7) <= maxPool4_CP_1841_elements(397);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	12 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	13 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_sample_start_
      -- CP-element group 8: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_request/$entry
      -- CP-element group 8: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_request/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_416_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(8), ack => addr_of_416_final_reg_req_0); -- 
    maxPool4_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(12) & maxPool4_CP_1841_elements(13);
      gj_maxPool4_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	38 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_update_start_
      -- CP-element group 9: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_complete/$entry
      -- CP-element group 9: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_complete/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_416_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(9), ack => addr_of_416_final_reg_req_1); -- 
    maxPool4_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(14) & maxPool4_CP_1841_elements(38);
      gj_maxPool4_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_final_index_sum_regn_Update/req
      -- CP-element group 10: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_final_index_sum_regn_update_start
      -- CP-element group 10: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_final_index_sum_regn_Update/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_415_index_offset_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(10), ack => array_obj_ref_415_index_offset_req_1); -- 
    maxPool4_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(12) & maxPool4_CP_1841_elements(13);
      gj_maxPool4_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	391 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	3 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_final_index_sum_regn_Sample/ack
      -- CP-element group 11: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_final_index_sum_regn_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_final_index_sum_regn_sample_complete
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_415_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_415_index_offset_ack_0, ack => maxPool4_CP_1841_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_offset_calculated
      -- CP-element group 12: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_root_address_calculated
      -- CP-element group 12: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_final_index_sum_regn_Update/ack
      -- CP-element group 12: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_final_index_sum_regn_Update/$exit
      -- CP-element group 12: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_base_plus_offset/$entry
      -- CP-element group 12: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_base_plus_offset/$exit
      -- CP-element group 12: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_base_plus_offset/sum_rename_req
      -- CP-element group 12: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_415_base_plus_offset/sum_rename_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_415_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_415_index_offset_ack_1, ack => maxPool4_CP_1841_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_sample_completed_
      -- CP-element group 13: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_request/$exit
      -- CP-element group 13: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_request/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_416_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_416_final_reg_ack_0, ack => maxPool4_CP_1841_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	9 
    -- CP-element group 14:  members (19) 
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_update_completed_
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_complete/ack
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_416_complete/$exit
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_base_address_resized
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_base_addr_resize/$entry
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_base_addr_resize/$exit
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_base_addr_resize/base_resize_req
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_base_addr_resize/base_resize_ack
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_base_plus_offset/$entry
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_base_plus_offset/$exit
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_base_plus_offset/sum_rename_req
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_base_plus_offset/sum_rename_ack
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_word_addrgen/$entry
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_word_addrgen/$exit
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_word_addrgen/root_register_req
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_word_addrgen/root_register_ack
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_base_address_calculated
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_word_address_calculated
      -- CP-element group 14: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_root_address_calculated
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_416_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_416_final_reg_ack_1, ack => maxPool4_CP_1841_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_request/req
      -- CP-element group 15: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_sample_start_
      -- CP-element group 15: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_request/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_423_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(15), ack => addr_of_423_final_reg_req_0); -- 
    maxPool4_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(19) & maxPool4_CP_1841_elements(20);
      gj_maxPool4_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	1 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	21 
    -- CP-element group 16: 	42 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_complete/$entry
      -- CP-element group 16: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_complete/req
      -- CP-element group 16: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_423_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(16), ack => addr_of_423_final_reg_req_1); -- 
    maxPool4_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(21) & maxPool4_CP_1841_elements(42);
      gj_maxPool4_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_final_index_sum_regn_Update/req
      -- CP-element group 17: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_final_index_sum_regn_Update/$entry
      -- CP-element group 17: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_final_index_sum_regn_update_start
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_422_index_offset_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(17), ack => array_obj_ref_422_index_offset_req_1); -- 
    maxPool4_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(19) & maxPool4_CP_1841_elements(20);
      gj_maxPool4_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	391 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	4 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_final_index_sum_regn_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_final_index_sum_regn_Sample/ack
      -- CP-element group 18: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_final_index_sum_regn_sample_complete
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_422_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_422_index_offset_ack_0, ack => maxPool4_CP_1841_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (8) 
      -- CP-element group 19: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_final_index_sum_regn_Update/$exit
      -- CP-element group 19: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_base_plus_offset/sum_rename_ack
      -- CP-element group 19: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_final_index_sum_regn_Update/ack
      -- CP-element group 19: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_base_plus_offset/$entry
      -- CP-element group 19: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_base_plus_offset/$exit
      -- CP-element group 19: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_offset_calculated
      -- CP-element group 19: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_422_root_address_calculated
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_422_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_422_index_offset_ack_1, ack => maxPool4_CP_1841_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_request/$exit
      -- CP-element group 20: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_request/ack
      -- CP-element group 20: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_423_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_423_final_reg_ack_0, ack => maxPool4_CP_1841_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	40 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21:  members (19) 
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_complete/$exit
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_complete/ack
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_423_update_completed_
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_base_address_calculated
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_word_address_calculated
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_root_address_calculated
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_base_address_resized
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_base_addr_resize/$entry
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_base_addr_resize/$exit
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_base_addr_resize/base_resize_req
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_base_plus_offset/$entry
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_base_plus_offset/$exit
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_word_addrgen/$entry
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_word_addrgen/$exit
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_word_addrgen/root_register_req
      -- CP-element group 21: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_423_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_423_final_reg_ack_1, ack => maxPool4_CP_1841_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	26 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	27 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_sample_start_
      -- CP-element group 22: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_request/$entry
      -- CP-element group 22: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_request/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_430_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(22), ack => addr_of_430_final_reg_req_0); -- 
    maxPool4_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(26) & maxPool4_CP_1841_elements(27);
      gj_maxPool4_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	1 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	28 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	28 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_complete/$entry
      -- CP-element group 23: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_update_start_
      -- CP-element group 23: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_complete/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_430_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(23), ack => addr_of_430_final_reg_req_1); -- 
    maxPool4_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(28) & maxPool4_CP_1841_elements(46);
      gj_maxPool4_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	1 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_final_index_sum_regn_update_start
      -- CP-element group 24: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_final_index_sum_regn_Update/$entry
      -- CP-element group 24: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_final_index_sum_regn_Update/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_429_index_offset_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(24), ack => array_obj_ref_429_index_offset_req_1); -- 
    maxPool4_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(26) & maxPool4_CP_1841_elements(27);
      gj_maxPool4_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	1 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	391 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	5 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_final_index_sum_regn_sample_complete
      -- CP-element group 25: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_final_index_sum_regn_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_429_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_429_index_offset_ack_0, ack => maxPool4_CP_1841_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	22 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (8) 
      -- CP-element group 26: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_root_address_calculated
      -- CP-element group 26: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_offset_calculated
      -- CP-element group 26: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_final_index_sum_regn_Update/$exit
      -- CP-element group 26: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_base_plus_offset/sum_rename_req
      -- CP-element group 26: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_final_index_sum_regn_Update/ack
      -- CP-element group 26: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_base_plus_offset/sum_rename_ack
      -- CP-element group 26: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_base_plus_offset/$entry
      -- CP-element group 26: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_429_base_plus_offset/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_429_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_429_index_offset_ack_1, ack => maxPool4_CP_1841_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: successors 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	24 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_sample_completed_
      -- CP-element group 27: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_request/ack
      -- CP-element group 27: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_request/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_430_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_430_final_reg_ack_0, ack => maxPool4_CP_1841_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	44 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	23 
    -- CP-element group 28:  members (19) 
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_update_completed_
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_complete/ack
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_430_complete/$exit
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_base_address_calculated
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_word_address_calculated
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_root_address_calculated
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_base_address_resized
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_base_addr_resize/$entry
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_base_addr_resize/$exit
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_base_addr_resize/base_resize_req
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_base_addr_resize/base_resize_ack
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_base_plus_offset/$entry
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_base_plus_offset/$exit
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_word_addrgen/$entry
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_word_addrgen/$exit
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_word_addrgen/root_register_req
      -- CP-element group 28: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_430_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_430_final_reg_ack_1, ack => maxPool4_CP_1841_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	33 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	34 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_sample_start_
      -- CP-element group 29: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_request/$entry
      -- CP-element group 29: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_request/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_437_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(29), ack => addr_of_437_final_reg_req_0); -- 
    maxPool4_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(33) & maxPool4_CP_1841_elements(34);
      gj_maxPool4_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	1 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	35 
    -- CP-element group 30: 	50 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	35 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_update_start_
      -- CP-element group 30: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_complete/$entry
      -- CP-element group 30: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_complete/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_437_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(30), ack => addr_of_437_final_reg_req_1); -- 
    maxPool4_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(35) & maxPool4_CP_1841_elements(50);
      gj_maxPool4_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	1 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	34 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_final_index_sum_regn_update_start
      -- CP-element group 31: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_final_index_sum_regn_Update/req
      -- CP-element group 31: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_final_index_sum_regn_Update/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_436_index_offset_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(31), ack => array_obj_ref_436_index_offset_req_1); -- 
    maxPool4_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(33) & maxPool4_CP_1841_elements(34);
      gj_maxPool4_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	1 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	391 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	6 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_final_index_sum_regn_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_final_index_sum_regn_Sample/ack
      -- CP-element group 32: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_final_index_sum_regn_sample_complete
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_436_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_436_index_offset_ack_0, ack => maxPool4_CP_1841_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	29 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (8) 
      -- CP-element group 33: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_offset_calculated
      -- CP-element group 33: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_final_index_sum_regn_Update/ack
      -- CP-element group 33: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_root_address_calculated
      -- CP-element group 33: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_final_index_sum_regn_Update/$exit
      -- CP-element group 33: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_base_plus_offset/$entry
      -- CP-element group 33: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_base_plus_offset/sum_rename_ack
      -- CP-element group 33: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_436_base_plus_offset/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_436_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_436_index_offset_ack_1, ack => maxPool4_CP_1841_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	31 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_sample_completed_
      -- CP-element group 34: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_request/$exit
      -- CP-element group 34: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_request/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_437_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_437_final_reg_ack_0, ack => maxPool4_CP_1841_elements(34)); -- 
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	30 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	48 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	30 
    -- CP-element group 35:  members (19) 
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_root_address_calculated
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_update_completed_
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_complete/ack
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_437_complete/$exit
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_base_address_calculated
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_word_address_calculated
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_base_address_resized
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_base_addr_resize/$entry
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_base_addr_resize/$exit
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_base_addr_resize/base_resize_req
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_base_addr_resize/base_resize_ack
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_base_plus_offset/$entry
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_base_plus_offset/$exit
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_word_addrgen/$entry
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_word_addrgen/$exit
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_word_addrgen/root_register_req
      -- CP-element group 35: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_437_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_437_final_reg_ack_1, ack => maxPool4_CP_1841_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Sample/word_access_start/word_0/$entry
      -- CP-element group 36: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Sample/word_access_start/word_0/rr
      -- CP-element group 36: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_sample_start_
      -- CP-element group 36: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Sample/$entry
      -- CP-element group 36: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Sample/word_access_start/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_441_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(36), ack => ptr_deref_441_load_0_req_0); -- 
    maxPool4_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(14) & maxPool4_CP_1841_elements(38);
      gj_maxPool4_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	54 
    -- CP-element group 37: 	58 
    -- CP-element group 37: 	62 
    -- CP-element group 37: 	66 
    -- CP-element group 37: 	70 
    -- CP-element group 37: 	74 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	82 
    -- CP-element group 37: 	86 
    -- CP-element group 37: 	90 
    -- CP-element group 37: 	94 
    -- CP-element group 37: 	98 
    -- CP-element group 37: 	102 
    -- CP-element group 37: 	106 
    -- CP-element group 37: 	110 
    -- CP-element group 37: 	114 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/$entry
      -- CP-element group 37: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/word_access_complete/$entry
      -- CP-element group 37: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/word_access_complete/word_0/cr
      -- CP-element group 37: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_441_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(37), ack => ptr_deref_441_load_0_req_1); -- 
    maxPool4_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(54) & maxPool4_CP_1841_elements(58) & maxPool4_CP_1841_elements(62) & maxPool4_CP_1841_elements(66) & maxPool4_CP_1841_elements(70) & maxPool4_CP_1841_elements(74) & maxPool4_CP_1841_elements(78) & maxPool4_CP_1841_elements(82) & maxPool4_CP_1841_elements(86) & maxPool4_CP_1841_elements(90) & maxPool4_CP_1841_elements(94) & maxPool4_CP_1841_elements(98) & maxPool4_CP_1841_elements(102) & maxPool4_CP_1841_elements(106) & maxPool4_CP_1841_elements(110) & maxPool4_CP_1841_elements(114);
      gj_maxPool4_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Sample/word_access_start/word_0/ra
      -- CP-element group 38: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Sample/$exit
      -- CP-element group 38: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Sample/word_access_start/$exit
      -- CP-element group 38: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_441_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_441_load_0_ack_0, ack => maxPool4_CP_1841_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	52 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	72 
    -- CP-element group 39: 	76 
    -- CP-element group 39: 	80 
    -- CP-element group 39: 	84 
    -- CP-element group 39: 	88 
    -- CP-element group 39: 	92 
    -- CP-element group 39: 	96 
    -- CP-element group 39: 	100 
    -- CP-element group 39: 	104 
    -- CP-element group 39: 	108 
    -- CP-element group 39: 	112 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/$exit
      -- CP-element group 39: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/word_access_complete/$exit
      -- CP-element group 39: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/ptr_deref_441_Merge/$entry
      -- CP-element group 39: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/ptr_deref_441_Merge/$exit
      -- CP-element group 39: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/ptr_deref_441_Merge/merge_req
      -- CP-element group 39: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_Update/ptr_deref_441_Merge/merge_ack
      -- CP-element group 39: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_441_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_441_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_441_load_0_ack_1, ack => maxPool4_CP_1841_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	21 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_sample_start_
      -- CP-element group 40: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Sample/$entry
      -- CP-element group 40: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Sample/word_access_start/$entry
      -- CP-element group 40: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Sample/word_access_start/word_0/$entry
      -- CP-element group 40: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_445_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(40), ack => ptr_deref_445_load_0_req_0); -- 
    maxPool4_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(21) & maxPool4_CP_1841_elements(42);
      gj_maxPool4_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	118 
    -- CP-element group 41: 	122 
    -- CP-element group 41: 	126 
    -- CP-element group 41: 	130 
    -- CP-element group 41: 	134 
    -- CP-element group 41: 	138 
    -- CP-element group 41: 	142 
    -- CP-element group 41: 	146 
    -- CP-element group 41: 	150 
    -- CP-element group 41: 	154 
    -- CP-element group 41: 	158 
    -- CP-element group 41: 	162 
    -- CP-element group 41: 	166 
    -- CP-element group 41: 	170 
    -- CP-element group 41: 	174 
    -- CP-element group 41: 	178 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_update_start_
      -- CP-element group 41: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/$entry
      -- CP-element group 41: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/word_access_complete/$entry
      -- CP-element group 41: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_445_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(41), ack => ptr_deref_445_load_0_req_1); -- 
    maxPool4_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(118) & maxPool4_CP_1841_elements(122) & maxPool4_CP_1841_elements(126) & maxPool4_CP_1841_elements(130) & maxPool4_CP_1841_elements(134) & maxPool4_CP_1841_elements(138) & maxPool4_CP_1841_elements(142) & maxPool4_CP_1841_elements(146) & maxPool4_CP_1841_elements(150) & maxPool4_CP_1841_elements(154) & maxPool4_CP_1841_elements(158) & maxPool4_CP_1841_elements(162) & maxPool4_CP_1841_elements(166) & maxPool4_CP_1841_elements(170) & maxPool4_CP_1841_elements(174) & maxPool4_CP_1841_elements(178);
      gj_maxPool4_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	16 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_sample_completed_
      -- CP-element group 42: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Sample/$exit
      -- CP-element group 42: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Sample/word_access_start/$exit
      -- CP-element group 42: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_445_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_445_load_0_ack_0, ack => maxPool4_CP_1841_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	116 
    -- CP-element group 43: 	120 
    -- CP-element group 43: 	124 
    -- CP-element group 43: 	128 
    -- CP-element group 43: 	132 
    -- CP-element group 43: 	136 
    -- CP-element group 43: 	140 
    -- CP-element group 43: 	144 
    -- CP-element group 43: 	148 
    -- CP-element group 43: 	152 
    -- CP-element group 43: 	156 
    -- CP-element group 43: 	160 
    -- CP-element group 43: 	164 
    -- CP-element group 43: 	168 
    -- CP-element group 43: 	172 
    -- CP-element group 43: 	176 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_update_completed_
      -- CP-element group 43: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/$exit
      -- CP-element group 43: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/word_access_complete/$exit
      -- CP-element group 43: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/ptr_deref_445_Merge/$entry
      -- CP-element group 43: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/ptr_deref_445_Merge/$exit
      -- CP-element group 43: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/ptr_deref_445_Merge/merge_req
      -- CP-element group 43: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_445_Update/ptr_deref_445_Merge/merge_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_445_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_445_load_0_ack_1, ack => maxPool4_CP_1841_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	28 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_sample_start_
      -- CP-element group 44: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Sample/$entry
      -- CP-element group 44: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Sample/word_access_start/$entry
      -- CP-element group 44: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_449_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(44), ack => ptr_deref_449_load_0_req_0); -- 
    maxPool4_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(28) & maxPool4_CP_1841_elements(46);
      gj_maxPool4_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: 	182 
    -- CP-element group 45: 	186 
    -- CP-element group 45: 	190 
    -- CP-element group 45: 	194 
    -- CP-element group 45: 	198 
    -- CP-element group 45: 	202 
    -- CP-element group 45: 	206 
    -- CP-element group 45: 	210 
    -- CP-element group 45: 	214 
    -- CP-element group 45: 	218 
    -- CP-element group 45: 	222 
    -- CP-element group 45: 	226 
    -- CP-element group 45: 	230 
    -- CP-element group 45: 	234 
    -- CP-element group 45: 	238 
    -- CP-element group 45: 	242 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_update_start_
      -- CP-element group 45: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/$entry
      -- CP-element group 45: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/word_access_complete/$entry
      -- CP-element group 45: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/word_access_complete/word_0/$entry
      -- CP-element group 45: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_449_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(45), ack => ptr_deref_449_load_0_req_1); -- 
    maxPool4_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(182) & maxPool4_CP_1841_elements(186) & maxPool4_CP_1841_elements(190) & maxPool4_CP_1841_elements(194) & maxPool4_CP_1841_elements(198) & maxPool4_CP_1841_elements(202) & maxPool4_CP_1841_elements(206) & maxPool4_CP_1841_elements(210) & maxPool4_CP_1841_elements(214) & maxPool4_CP_1841_elements(218) & maxPool4_CP_1841_elements(222) & maxPool4_CP_1841_elements(226) & maxPool4_CP_1841_elements(230) & maxPool4_CP_1841_elements(234) & maxPool4_CP_1841_elements(238) & maxPool4_CP_1841_elements(242);
      gj_maxPool4_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_sample_completed_
      -- CP-element group 46: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Sample/$exit
      -- CP-element group 46: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Sample/word_access_start/$exit
      -- CP-element group 46: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_449_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_449_load_0_ack_0, ack => maxPool4_CP_1841_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	180 
    -- CP-element group 47: 	184 
    -- CP-element group 47: 	188 
    -- CP-element group 47: 	192 
    -- CP-element group 47: 	196 
    -- CP-element group 47: 	200 
    -- CP-element group 47: 	204 
    -- CP-element group 47: 	208 
    -- CP-element group 47: 	212 
    -- CP-element group 47: 	216 
    -- CP-element group 47: 	220 
    -- CP-element group 47: 	224 
    -- CP-element group 47: 	228 
    -- CP-element group 47: 	232 
    -- CP-element group 47: 	236 
    -- CP-element group 47: 	240 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_update_completed_
      -- CP-element group 47: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/$exit
      -- CP-element group 47: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/word_access_complete/$exit
      -- CP-element group 47: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/word_access_complete/word_0/ca
      -- CP-element group 47: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/ptr_deref_449_Merge/$entry
      -- CP-element group 47: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/ptr_deref_449_Merge/$exit
      -- CP-element group 47: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/ptr_deref_449_Merge/merge_req
      -- CP-element group 47: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_449_Update/ptr_deref_449_Merge/merge_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_449_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_449_load_0_ack_1, ack => maxPool4_CP_1841_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	35 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_sample_start_
      -- CP-element group 48: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Sample/$entry
      -- CP-element group 48: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Sample/word_access_start/$entry
      -- CP-element group 48: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_453_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(48), ack => ptr_deref_453_load_0_req_0); -- 
    maxPool4_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(35) & maxPool4_CP_1841_elements(50);
      gj_maxPool4_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: 	246 
    -- CP-element group 49: 	250 
    -- CP-element group 49: 	254 
    -- CP-element group 49: 	258 
    -- CP-element group 49: 	262 
    -- CP-element group 49: 	266 
    -- CP-element group 49: 	270 
    -- CP-element group 49: 	274 
    -- CP-element group 49: 	278 
    -- CP-element group 49: 	282 
    -- CP-element group 49: 	286 
    -- CP-element group 49: 	290 
    -- CP-element group 49: 	294 
    -- CP-element group 49: 	298 
    -- CP-element group 49: 	302 
    -- CP-element group 49: 	306 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_update_start_
      -- CP-element group 49: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/$entry
      -- CP-element group 49: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/word_access_complete/$entry
      -- CP-element group 49: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/word_access_complete/word_0/$entry
      -- CP-element group 49: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_453_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(49), ack => ptr_deref_453_load_0_req_1); -- 
    maxPool4_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(246) & maxPool4_CP_1841_elements(250) & maxPool4_CP_1841_elements(254) & maxPool4_CP_1841_elements(258) & maxPool4_CP_1841_elements(262) & maxPool4_CP_1841_elements(266) & maxPool4_CP_1841_elements(270) & maxPool4_CP_1841_elements(274) & maxPool4_CP_1841_elements(278) & maxPool4_CP_1841_elements(282) & maxPool4_CP_1841_elements(286) & maxPool4_CP_1841_elements(290) & maxPool4_CP_1841_elements(294) & maxPool4_CP_1841_elements(298) & maxPool4_CP_1841_elements(302) & maxPool4_CP_1841_elements(306);
      gj_maxPool4_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	30 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_sample_completed_
      -- CP-element group 50: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Sample/$exit
      -- CP-element group 50: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Sample/word_access_start/$exit
      -- CP-element group 50: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_453_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_453_load_0_ack_0, ack => maxPool4_CP_1841_elements(50)); -- 
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	244 
    -- CP-element group 51: 	248 
    -- CP-element group 51: 	252 
    -- CP-element group 51: 	256 
    -- CP-element group 51: 	260 
    -- CP-element group 51: 	264 
    -- CP-element group 51: 	268 
    -- CP-element group 51: 	272 
    -- CP-element group 51: 	276 
    -- CP-element group 51: 	280 
    -- CP-element group 51: 	284 
    -- CP-element group 51: 	288 
    -- CP-element group 51: 	292 
    -- CP-element group 51: 	296 
    -- CP-element group 51: 	300 
    -- CP-element group 51: 	304 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_update_completed_
      -- CP-element group 51: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/$exit
      -- CP-element group 51: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/word_access_complete/$exit
      -- CP-element group 51: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/word_access_complete/word_0/ca
      -- CP-element group 51: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/ptr_deref_453_Merge/$entry
      -- CP-element group 51: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/ptr_deref_453_Merge/$exit
      -- CP-element group 51: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/ptr_deref_453_Merge/merge_req
      -- CP-element group 51: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_453_Update/ptr_deref_453_Merge/merge_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_453_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_453_load_0_ack_1, ack => maxPool4_CP_1841_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	39 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_sample_start_
      -- CP-element group 52: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_Sample/$entry
      -- CP-element group 52: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_457_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(52), ack => slice_457_inst_req_0); -- 
    maxPool4_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(54);
      gj_maxPool4_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	321 
    -- CP-element group 53: 	386 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_update_start_
      -- CP-element group 53: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_Update/$entry
      -- CP-element group 53: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_457_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(53), ack => slice_457_inst_req_1); -- 
    maxPool4_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(55) & maxPool4_CP_1841_elements(321) & maxPool4_CP_1841_elements(386);
      gj_maxPool4_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	37 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_sample_completed_
      -- CP-element group 54: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_Sample/$exit
      -- CP-element group 54: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_457_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_457_inst_ack_0, ack => maxPool4_CP_1841_elements(54)); -- 
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	319 
    -- CP-element group 55: 	384 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_update_completed_
      -- CP-element group 55: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_Update/$exit
      -- CP-element group 55: 	 assign_stmt_417_to_assign_stmt_1457/slice_457_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_457_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_457_inst_ack_1, ack => maxPool4_CP_1841_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_sample_start_
      -- CP-element group 56: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_Sample/$entry
      -- CP-element group 56: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_461_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(56), ack => slice_461_inst_req_0); -- 
    maxPool4_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(58);
      gj_maxPool4_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	321 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_update_start_
      -- CP-element group 57: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_Update/$entry
      -- CP-element group 57: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_461_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(57), ack => slice_461_inst_req_1); -- 
    maxPool4_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(59) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	37 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_sample_completed_
      -- CP-element group 58: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_Sample/$exit
      -- CP-element group 58: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_461_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_461_inst_ack_0, ack => maxPool4_CP_1841_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	319 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_update_completed_
      -- CP-element group 59: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_Update/$exit
      -- CP-element group 59: 	 assign_stmt_417_to_assign_stmt_1457/slice_461_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_461_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_461_inst_ack_1, ack => maxPool4_CP_1841_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_sample_start_
      -- CP-element group 60: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_Sample/$entry
      -- CP-element group 60: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_465_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(60), ack => slice_465_inst_req_0); -- 
    maxPool4_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(62);
      gj_maxPool4_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	321 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_update_start_
      -- CP-element group 61: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_Update/$entry
      -- CP-element group 61: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_465_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(61), ack => slice_465_inst_req_1); -- 
    maxPool4_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(63) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	37 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_sample_completed_
      -- CP-element group 62: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_Sample/$exit
      -- CP-element group 62: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_465_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_465_inst_ack_0, ack => maxPool4_CP_1841_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	319 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_update_completed_
      -- CP-element group 63: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_Update/$exit
      -- CP-element group 63: 	 assign_stmt_417_to_assign_stmt_1457/slice_465_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_465_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_465_inst_ack_1, ack => maxPool4_CP_1841_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_sample_start_
      -- CP-element group 64: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_Sample/$entry
      -- CP-element group 64: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_469_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(64), ack => slice_469_inst_req_0); -- 
    maxPool4_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(66);
      gj_maxPool4_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	321 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_update_start_
      -- CP-element group 65: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_Update/$entry
      -- CP-element group 65: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_469_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(65), ack => slice_469_inst_req_1); -- 
    maxPool4_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(67) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	37 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_sample_completed_
      -- CP-element group 66: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_Sample/$exit
      -- CP-element group 66: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_469_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_469_inst_ack_0, ack => maxPool4_CP_1841_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	319 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_update_completed_
      -- CP-element group 67: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_Update/$exit
      -- CP-element group 67: 	 assign_stmt_417_to_assign_stmt_1457/slice_469_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_469_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_469_inst_ack_1, ack => maxPool4_CP_1841_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_sample_start_
      -- CP-element group 68: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_Sample/$entry
      -- CP-element group 68: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_473_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(68), ack => slice_473_inst_req_0); -- 
    maxPool4_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(70);
      gj_maxPool4_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: 	340 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_update_start_
      -- CP-element group 69: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_Update/$entry
      -- CP-element group 69: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_473_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(69), ack => slice_473_inst_req_1); -- 
    maxPool4_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(71) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	37 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_sample_completed_
      -- CP-element group 70: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_Sample/$exit
      -- CP-element group 70: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_473_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_473_inst_ack_0, ack => maxPool4_CP_1841_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	338 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_update_completed_
      -- CP-element group 71: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_Update/$exit
      -- CP-element group 71: 	 assign_stmt_417_to_assign_stmt_1457/slice_473_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_473_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_473_inst_ack_1, ack => maxPool4_CP_1841_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	39 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_sample_start_
      -- CP-element group 72: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_Sample/$entry
      -- CP-element group 72: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_477_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(72), ack => slice_477_inst_req_0); -- 
    maxPool4_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(74);
      gj_maxPool4_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: 	340 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_update_start_
      -- CP-element group 73: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_Update/$entry
      -- CP-element group 73: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_477_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(73), ack => slice_477_inst_req_1); -- 
    maxPool4_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(75) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	37 
    -- CP-element group 74: 	72 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_sample_completed_
      -- CP-element group 74: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_Sample/$exit
      -- CP-element group 74: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_477_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_477_inst_ack_0, ack => maxPool4_CP_1841_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	338 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_update_completed_
      -- CP-element group 75: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_Update/$exit
      -- CP-element group 75: 	 assign_stmt_417_to_assign_stmt_1457/slice_477_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_477_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_477_inst_ack_1, ack => maxPool4_CP_1841_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	39 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_sample_start_
      -- CP-element group 76: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_Sample/$entry
      -- CP-element group 76: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_481_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(76), ack => slice_481_inst_req_0); -- 
    maxPool4_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(78);
      gj_maxPool4_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	340 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_update_start_
      -- CP-element group 77: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_Update/$entry
      -- CP-element group 77: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_481_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(77), ack => slice_481_inst_req_1); -- 
    maxPool4_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(79) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_sample_completed_
      -- CP-element group 78: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_Sample/$exit
      -- CP-element group 78: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_481_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_481_inst_ack_0, ack => maxPool4_CP_1841_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	338 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_update_completed_
      -- CP-element group 79: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_Update/$exit
      -- CP-element group 79: 	 assign_stmt_417_to_assign_stmt_1457/slice_481_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_481_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_481_inst_ack_1, ack => maxPool4_CP_1841_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	39 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_sample_start_
      -- CP-element group 80: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_Sample/$entry
      -- CP-element group 80: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_485_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(80), ack => slice_485_inst_req_0); -- 
    maxPool4_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(82);
      gj_maxPool4_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: 	340 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_update_start_
      -- CP-element group 81: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_Update/$entry
      -- CP-element group 81: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_485_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(81), ack => slice_485_inst_req_1); -- 
    maxPool4_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(83) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	37 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_sample_completed_
      -- CP-element group 82: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_Sample/$exit
      -- CP-element group 82: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_485_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_485_inst_ack_0, ack => maxPool4_CP_1841_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	338 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_update_completed_
      -- CP-element group 83: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_Update/$exit
      -- CP-element group 83: 	 assign_stmt_417_to_assign_stmt_1457/slice_485_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_485_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_485_inst_ack_1, ack => maxPool4_CP_1841_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	39 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_sample_start_
      -- CP-element group 84: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_Sample/$entry
      -- CP-element group 84: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_489_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(84), ack => slice_489_inst_req_0); -- 
    maxPool4_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(86);
      gj_maxPool4_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: 	359 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_update_start_
      -- CP-element group 85: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_Update/$entry
      -- CP-element group 85: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_489_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(85), ack => slice_489_inst_req_1); -- 
    maxPool4_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(87) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	37 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_sample_completed_
      -- CP-element group 86: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_Sample/$exit
      -- CP-element group 86: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_489_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_489_inst_ack_0, ack => maxPool4_CP_1841_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	357 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_update_completed_
      -- CP-element group 87: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_Update/$exit
      -- CP-element group 87: 	 assign_stmt_417_to_assign_stmt_1457/slice_489_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_489_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_489_inst_ack_1, ack => maxPool4_CP_1841_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	39 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_sample_start_
      -- CP-element group 88: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_Sample/$entry
      -- CP-element group 88: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_493_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(88), ack => slice_493_inst_req_0); -- 
    maxPool4_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(90);
      gj_maxPool4_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: 	359 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_update_start_
      -- CP-element group 89: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_Update/$entry
      -- CP-element group 89: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_493_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(89), ack => slice_493_inst_req_1); -- 
    maxPool4_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(91) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	37 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_sample_completed_
      -- CP-element group 90: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_Sample/$exit
      -- CP-element group 90: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_493_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_493_inst_ack_0, ack => maxPool4_CP_1841_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	357 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_update_completed_
      -- CP-element group 91: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_Update/$exit
      -- CP-element group 91: 	 assign_stmt_417_to_assign_stmt_1457/slice_493_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_493_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_493_inst_ack_1, ack => maxPool4_CP_1841_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	39 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_sample_start_
      -- CP-element group 92: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_Sample/$entry
      -- CP-element group 92: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_497_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(92), ack => slice_497_inst_req_0); -- 
    maxPool4_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(94);
      gj_maxPool4_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: 	359 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_update_start_
      -- CP-element group 93: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_Update/$entry
      -- CP-element group 93: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_497_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(93), ack => slice_497_inst_req_1); -- 
    maxPool4_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(95) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	37 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_sample_completed_
      -- CP-element group 94: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_Sample/$exit
      -- CP-element group 94: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_497_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_497_inst_ack_0, ack => maxPool4_CP_1841_elements(94)); -- 
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	357 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_update_completed_
      -- CP-element group 95: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_Update/$exit
      -- CP-element group 95: 	 assign_stmt_417_to_assign_stmt_1457/slice_497_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_497_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_497_inst_ack_1, ack => maxPool4_CP_1841_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	39 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_sample_start_
      -- CP-element group 96: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_Sample/$entry
      -- CP-element group 96: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_501_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(96), ack => slice_501_inst_req_0); -- 
    maxPool4_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(98);
      gj_maxPool4_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	359 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_update_start_
      -- CP-element group 97: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_Update/$entry
      -- CP-element group 97: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_501_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(97), ack => slice_501_inst_req_1); -- 
    maxPool4_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(99) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	37 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_sample_completed_
      -- CP-element group 98: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_Sample/$exit
      -- CP-element group 98: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_501_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_501_inst_ack_0, ack => maxPool4_CP_1841_elements(98)); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	357 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_update_completed_
      -- CP-element group 99: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_Update/$exit
      -- CP-element group 99: 	 assign_stmt_417_to_assign_stmt_1457/slice_501_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_501_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_501_inst_ack_1, ack => maxPool4_CP_1841_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	39 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_sample_start_
      -- CP-element group 100: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_Sample/$entry
      -- CP-element group 100: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(100) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_505_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(100), ack => slice_505_inst_req_0); -- 
    maxPool4_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(102);
      gj_maxPool4_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: 	378 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_update_start_
      -- CP-element group 101: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_Update/$entry
      -- CP-element group 101: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_505_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(101), ack => slice_505_inst_req_1); -- 
    maxPool4_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(103) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	37 
    -- CP-element group 102: 	100 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_sample_completed_
      -- CP-element group 102: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_Sample/$exit
      -- CP-element group 102: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_505_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_505_inst_ack_0, ack => maxPool4_CP_1841_elements(102)); -- 
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	376 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_update_completed_
      -- CP-element group 103: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_Update/$exit
      -- CP-element group 103: 	 assign_stmt_417_to_assign_stmt_1457/slice_505_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(103) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_505_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_505_inst_ack_1, ack => maxPool4_CP_1841_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	39 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_sample_start_
      -- CP-element group 104: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_Sample/$entry
      -- CP-element group 104: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_509_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(104), ack => slice_509_inst_req_0); -- 
    maxPool4_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(106);
      gj_maxPool4_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	378 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_update_start_
      -- CP-element group 105: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_Update/$entry
      -- CP-element group 105: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_509_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(105), ack => slice_509_inst_req_1); -- 
    maxPool4_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(107) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	37 
    -- CP-element group 106: 	104 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_sample_completed_
      -- CP-element group 106: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_Sample/$exit
      -- CP-element group 106: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_509_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_509_inst_ack_0, ack => maxPool4_CP_1841_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	376 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_update_completed_
      -- CP-element group 107: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_Update/$exit
      -- CP-element group 107: 	 assign_stmt_417_to_assign_stmt_1457/slice_509_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_509_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_509_inst_ack_1, ack => maxPool4_CP_1841_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	39 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_sample_start_
      -- CP-element group 108: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_Sample/$entry
      -- CP-element group 108: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_513_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(108), ack => slice_513_inst_req_0); -- 
    maxPool4_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(110);
      gj_maxPool4_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	378 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_update_start_
      -- CP-element group 109: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_Update/$entry
      -- CP-element group 109: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_513_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(109), ack => slice_513_inst_req_1); -- 
    maxPool4_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(111) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	37 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_sample_completed_
      -- CP-element group 110: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_Sample/$exit
      -- CP-element group 110: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_513_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_513_inst_ack_0, ack => maxPool4_CP_1841_elements(110)); -- 
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	376 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_update_completed_
      -- CP-element group 111: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_Update/$exit
      -- CP-element group 111: 	 assign_stmt_417_to_assign_stmt_1457/slice_513_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_513_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_513_inst_ack_1, ack => maxPool4_CP_1841_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	39 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_sample_start_
      -- CP-element group 112: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_Sample/$entry
      -- CP-element group 112: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_517_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(112), ack => slice_517_inst_req_0); -- 
    maxPool4_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(39) & maxPool4_CP_1841_elements(114);
      gj_maxPool4_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: 	378 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_update_start_
      -- CP-element group 113: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_Update/$entry
      -- CP-element group 113: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_517_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(113), ack => slice_517_inst_req_1); -- 
    maxPool4_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(115) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	37 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_sample_completed_
      -- CP-element group 114: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_Sample/$exit
      -- CP-element group 114: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_517_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_517_inst_ack_0, ack => maxPool4_CP_1841_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	376 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_update_completed_
      -- CP-element group 115: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_Update/$exit
      -- CP-element group 115: 	 assign_stmt_417_to_assign_stmt_1457/slice_517_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_517_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_517_inst_ack_1, ack => maxPool4_CP_1841_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	43 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_sample_start_
      -- CP-element group 116: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_Sample/$entry
      -- CP-element group 116: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_521_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(116), ack => slice_521_inst_req_0); -- 
    maxPool4_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(118);
      gj_maxPool4_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: 	321 
    -- CP-element group 117: 	386 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_update_start_
      -- CP-element group 117: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_Update/$entry
      -- CP-element group 117: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_521_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(117), ack => slice_521_inst_req_1); -- 
    maxPool4_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(119) & maxPool4_CP_1841_elements(321) & maxPool4_CP_1841_elements(386);
      gj_maxPool4_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	41 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_sample_completed_
      -- CP-element group 118: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_Sample/$exit
      -- CP-element group 118: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(118) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_521_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_521_inst_ack_0, ack => maxPool4_CP_1841_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	319 
    -- CP-element group 119: 	384 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	117 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_update_completed_
      -- CP-element group 119: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_Update/$exit
      -- CP-element group 119: 	 assign_stmt_417_to_assign_stmt_1457/slice_521_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_521_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_521_inst_ack_1, ack => maxPool4_CP_1841_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	43 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_sample_start_
      -- CP-element group 120: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_Sample/$entry
      -- CP-element group 120: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_525_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(120), ack => slice_525_inst_req_0); -- 
    maxPool4_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(122);
      gj_maxPool4_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	321 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_update_start_
      -- CP-element group 121: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_Update/$entry
      -- CP-element group 121: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_525_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(121), ack => slice_525_inst_req_1); -- 
    maxPool4_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(123) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	41 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_sample_completed_
      -- CP-element group 122: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_Sample/$exit
      -- CP-element group 122: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(122) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_525_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_525_inst_ack_0, ack => maxPool4_CP_1841_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	319 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	121 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_update_completed_
      -- CP-element group 123: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_Update/$exit
      -- CP-element group 123: 	 assign_stmt_417_to_assign_stmt_1457/slice_525_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_525_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_525_inst_ack_1, ack => maxPool4_CP_1841_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	43 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_sample_start_
      -- CP-element group 124: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_Sample/$entry
      -- CP-element group 124: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_529_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(124), ack => slice_529_inst_req_0); -- 
    maxPool4_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(126);
      gj_maxPool4_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: 	321 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_update_start_
      -- CP-element group 125: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_Update/$entry
      -- CP-element group 125: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_529_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(125), ack => slice_529_inst_req_1); -- 
    maxPool4_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(127) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	41 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_sample_completed_
      -- CP-element group 126: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_Sample/$exit
      -- CP-element group 126: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_529_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_529_inst_ack_0, ack => maxPool4_CP_1841_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	319 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_update_completed_
      -- CP-element group 127: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_Update/$exit
      -- CP-element group 127: 	 assign_stmt_417_to_assign_stmt_1457/slice_529_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_529_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_529_inst_ack_1, ack => maxPool4_CP_1841_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	43 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_sample_start_
      -- CP-element group 128: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_Sample/$entry
      -- CP-element group 128: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_533_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(128), ack => slice_533_inst_req_0); -- 
    maxPool4_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(130);
      gj_maxPool4_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: 	321 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_update_start_
      -- CP-element group 129: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_Update/$entry
      -- CP-element group 129: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_533_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(129), ack => slice_533_inst_req_1); -- 
    maxPool4_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(131) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	41 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_sample_completed_
      -- CP-element group 130: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_Sample/$exit
      -- CP-element group 130: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_533_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_533_inst_ack_0, ack => maxPool4_CP_1841_elements(130)); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	319 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_update_completed_
      -- CP-element group 131: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_Update/$exit
      -- CP-element group 131: 	 assign_stmt_417_to_assign_stmt_1457/slice_533_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(131) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_533_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_533_inst_ack_1, ack => maxPool4_CP_1841_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	43 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_Sample/rr
      -- CP-element group 132: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_Sample/$entry
      -- CP-element group 132: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(132) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_537_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(132), ack => slice_537_inst_req_0); -- 
    maxPool4_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(134);
      gj_maxPool4_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: 	340 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_Update/cr
      -- CP-element group 133: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_Update/$entry
      -- CP-element group 133: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(133) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_537_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(133), ack => slice_537_inst_req_1); -- 
    maxPool4_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(135) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	41 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_Sample/ra
      -- CP-element group 134: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_Sample/$exit
      -- CP-element group 134: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(134) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_537_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_537_inst_ack_0, ack => maxPool4_CP_1841_elements(134)); -- 
    -- CP-element group 135:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	338 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_Update/ca
      -- CP-element group 135: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_Update/$exit
      -- CP-element group 135: 	 assign_stmt_417_to_assign_stmt_1457/slice_537_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(135) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_537_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_537_inst_ack_1, ack => maxPool4_CP_1841_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	43 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_Sample/$entry
      -- CP-element group 136: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_Sample/rr
      -- CP-element group 136: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(136) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_541_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(136), ack => slice_541_inst_req_0); -- 
    maxPool4_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(138);
      gj_maxPool4_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: 	340 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_Update/cr
      -- CP-element group 137: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_Update/$entry
      -- CP-element group 137: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(137) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_541_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(137), ack => slice_541_inst_req_1); -- 
    maxPool4_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(139) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	41 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_Sample/$exit
      -- CP-element group 138: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_Sample/ra
      -- CP-element group 138: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_541_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_541_inst_ack_0, ack => maxPool4_CP_1841_elements(138)); -- 
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	338 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_Update/ca
      -- CP-element group 139: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_update_completed_
      -- CP-element group 139: 	 assign_stmt_417_to_assign_stmt_1457/slice_541_Update/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(139) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_541_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_541_inst_ack_1, ack => maxPool4_CP_1841_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	43 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_Sample/rr
      -- CP-element group 140: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_sample_start_
      -- CP-element group 140: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_Sample/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_545_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(140), ack => slice_545_inst_req_0); -- 
    maxPool4_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(142);
      gj_maxPool4_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: 	340 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_update_start_
      -- CP-element group 141: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_Update/$entry
      -- CP-element group 141: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(141) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_545_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(141), ack => slice_545_inst_req_1); -- 
    maxPool4_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(143) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	41 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_Sample/ra
      -- CP-element group 142: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_sample_completed_
      -- CP-element group 142: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_Sample/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(142) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_545_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_545_inst_ack_0, ack => maxPool4_CP_1841_elements(142)); -- 
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	338 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_Update/ca
      -- CP-element group 143: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_Update/$exit
      -- CP-element group 143: 	 assign_stmt_417_to_assign_stmt_1457/slice_545_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(143) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_545_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_545_inst_ack_1, ack => maxPool4_CP_1841_elements(143)); -- 
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	43 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_Sample/rr
      -- CP-element group 144: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_Sample/$entry
      -- CP-element group 144: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(144) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_549_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(144), ack => slice_549_inst_req_0); -- 
    maxPool4_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(146);
      gj_maxPool4_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: 	340 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_Update/cr
      -- CP-element group 145: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_Update/$entry
      -- CP-element group 145: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(145) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_549_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(145), ack => slice_549_inst_req_1); -- 
    maxPool4_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(147) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	41 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_Sample/ra
      -- CP-element group 146: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_Sample/$exit
      -- CP-element group 146: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(146) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_549_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_549_inst_ack_0, ack => maxPool4_CP_1841_elements(146)); -- 
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	338 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_Update/ca
      -- CP-element group 147: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_Update/$exit
      -- CP-element group 147: 	 assign_stmt_417_to_assign_stmt_1457/slice_549_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(147) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_549_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_549_inst_ack_1, ack => maxPool4_CP_1841_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	43 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_Sample/rr
      -- CP-element group 148: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_Sample/$entry
      -- CP-element group 148: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(148) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_553_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(148), ack => slice_553_inst_req_0); -- 
    maxPool4_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(150);
      gj_maxPool4_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: 	359 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_update_start_
      -- CP-element group 149: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_Update/$entry
      -- CP-element group 149: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(149) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_553_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(149), ack => slice_553_inst_req_1); -- 
    maxPool4_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(151) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	41 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_Sample/$exit
      -- CP-element group 150: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_sample_completed_
      -- CP-element group 150: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(150) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_553_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_553_inst_ack_0, ack => maxPool4_CP_1841_elements(150)); -- 
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	357 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_update_completed_
      -- CP-element group 151: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_Update/$exit
      -- CP-element group 151: 	 assign_stmt_417_to_assign_stmt_1457/slice_553_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(151) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_553_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_553_inst_ack_1, ack => maxPool4_CP_1841_elements(151)); -- 
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	43 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_sample_start_
      -- CP-element group 152: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_Sample/rr
      -- CP-element group 152: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_Sample/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(152) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_557_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(152), ack => slice_557_inst_req_0); -- 
    maxPool4_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(154);
      gj_maxPool4_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: 	359 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_update_start_
      -- CP-element group 153: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_Update/cr
      -- CP-element group 153: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_Update/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(153) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_557_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(153), ack => slice_557_inst_req_1); -- 
    maxPool4_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(155) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	41 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_sample_completed_
      -- CP-element group 154: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_Sample/ra
      -- CP-element group 154: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_Sample/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(154) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_557_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_557_inst_ack_0, ack => maxPool4_CP_1841_elements(154)); -- 
    -- CP-element group 155:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	357 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_update_completed_
      -- CP-element group 155: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_Update/ca
      -- CP-element group 155: 	 assign_stmt_417_to_assign_stmt_1457/slice_557_Update/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(155) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_557_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_557_inst_ack_1, ack => maxPool4_CP_1841_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	43 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_Sample/rr
      -- CP-element group 156: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_Sample/$entry
      -- CP-element group 156: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_561_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(156), ack => slice_561_inst_req_0); -- 
    maxPool4_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(158);
      gj_maxPool4_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: 	359 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_Update/cr
      -- CP-element group 157: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_Update/$entry
      -- CP-element group 157: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_561_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(157), ack => slice_561_inst_req_1); -- 
    maxPool4_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(159) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	41 
    -- CP-element group 158: 	156 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_Sample/ra
      -- CP-element group 158: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_Sample/$exit
      -- CP-element group 158: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(158) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_561_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_561_inst_ack_0, ack => maxPool4_CP_1841_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	357 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_Update/$exit
      -- CP-element group 159: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_update_completed_
      -- CP-element group 159: 	 assign_stmt_417_to_assign_stmt_1457/slice_561_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_561_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_561_inst_ack_1, ack => maxPool4_CP_1841_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	43 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_Sample/rr
      -- CP-element group 160: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_Sample/$entry
      -- CP-element group 160: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(160) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_565_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(160), ack => slice_565_inst_req_0); -- 
    maxPool4_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(162);
      gj_maxPool4_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: 	359 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_Update/cr
      -- CP-element group 161: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_Update/$entry
      -- CP-element group 161: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(161) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_565_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(161), ack => slice_565_inst_req_1); -- 
    maxPool4_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(163) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	41 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_Sample/ra
      -- CP-element group 162: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_Sample/$exit
      -- CP-element group 162: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_565_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_565_inst_ack_0, ack => maxPool4_CP_1841_elements(162)); -- 
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	357 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_Update/ca
      -- CP-element group 163: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_Update/$exit
      -- CP-element group 163: 	 assign_stmt_417_to_assign_stmt_1457/slice_565_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_565_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_565_inst_ack_1, ack => maxPool4_CP_1841_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	43 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_Sample/rr
      -- CP-element group 164: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_Sample/$entry
      -- CP-element group 164: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(164) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_569_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(164), ack => slice_569_inst_req_0); -- 
    maxPool4_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(166);
      gj_maxPool4_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: 	378 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_Update/cr
      -- CP-element group 165: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_Update/$entry
      -- CP-element group 165: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_569_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(165), ack => slice_569_inst_req_1); -- 
    maxPool4_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(167) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	41 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_Sample/ra
      -- CP-element group 166: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_Sample/$exit
      -- CP-element group 166: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(166) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_569_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_569_inst_ack_0, ack => maxPool4_CP_1841_elements(166)); -- 
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	376 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	165 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_Update/ca
      -- CP-element group 167: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_Update/$exit
      -- CP-element group 167: 	 assign_stmt_417_to_assign_stmt_1457/slice_569_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_569_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_569_inst_ack_1, ack => maxPool4_CP_1841_elements(167)); -- 
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	43 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_Sample/rr
      -- CP-element group 168: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_Sample/$entry
      -- CP-element group 168: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(168)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(168)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(168) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_573_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(168), ack => slice_573_inst_req_0); -- 
    maxPool4_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(170);
      gj_maxPool4_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: 	378 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_Update/cr
      -- CP-element group 169: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_Update/$entry
      -- CP-element group 169: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(169)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(169)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(169) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_573_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(169), ack => slice_573_inst_req_1); -- 
    maxPool4_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(171) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	41 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_Sample/ra
      -- CP-element group 170: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_Sample/$exit
      -- CP-element group 170: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(170)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(170)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(170) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_573_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_573_inst_ack_0, ack => maxPool4_CP_1841_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	376 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_Update/ca
      -- CP-element group 171: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_Update/$exit
      -- CP-element group 171: 	 assign_stmt_417_to_assign_stmt_1457/slice_573_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(171)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(171)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(171) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_573_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_573_inst_ack_1, ack => maxPool4_CP_1841_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	43 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_Sample/rr
      -- CP-element group 172: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_Sample/$entry
      -- CP-element group 172: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(172)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(172)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(172) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_577_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(172), ack => slice_577_inst_req_0); -- 
    maxPool4_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(174);
      gj_maxPool4_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: 	378 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_Update/cr
      -- CP-element group 173: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_Update/$entry
      -- CP-element group 173: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(173)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(173)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(173) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_577_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(173), ack => slice_577_inst_req_1); -- 
    maxPool4_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(175) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	41 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_Sample/ra
      -- CP-element group 174: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_Sample/$exit
      -- CP-element group 174: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(174)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(174)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(174) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_577_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_577_inst_ack_0, ack => maxPool4_CP_1841_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	376 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_Update/ca
      -- CP-element group 175: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_Update/$exit
      -- CP-element group 175: 	 assign_stmt_417_to_assign_stmt_1457/slice_577_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(175)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(175)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(175) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_577_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_577_inst_ack_1, ack => maxPool4_CP_1841_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	43 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_Sample/rr
      -- CP-element group 176: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_Sample/$entry
      -- CP-element group 176: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(176)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(176)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(176) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_581_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(176), ack => slice_581_inst_req_0); -- 
    maxPool4_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(43) & maxPool4_CP_1841_elements(178);
      gj_maxPool4_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: 	378 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_update_start_
      -- CP-element group 177: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_Update/cr
      -- CP-element group 177: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_Update/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(177)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(177)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(177) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_581_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(177), ack => slice_581_inst_req_1); -- 
    maxPool4_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(179) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	41 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_Sample/ra
      -- CP-element group 178: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_Sample/$exit
      -- CP-element group 178: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(178)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(178)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(178) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_581_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_581_inst_ack_0, ack => maxPool4_CP_1841_elements(178)); -- 
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	376 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_Update/ca
      -- CP-element group 179: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_Update/$exit
      -- CP-element group 179: 	 assign_stmt_417_to_assign_stmt_1457/slice_581_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(179)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(179)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(179) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_581_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_581_inst_ack_1, ack => maxPool4_CP_1841_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	47 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_Sample/$entry
      -- CP-element group 180: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_sample_start_
      -- CP-element group 180: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(180)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(180)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(180) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_585_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(180), ack => slice_585_inst_req_0); -- 
    maxPool4_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(182);
      gj_maxPool4_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: 	321 
    -- CP-element group 181: 	386 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_Update/$entry
      -- CP-element group 181: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_update_start_
      -- CP-element group 181: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(181)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(181)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(181) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_585_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(181), ack => slice_585_inst_req_1); -- 
    maxPool4_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(183) & maxPool4_CP_1841_elements(321) & maxPool4_CP_1841_elements(386);
      gj_maxPool4_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	45 
    -- CP-element group 182: 	180 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_Sample/ra
      -- CP-element group 182: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_Sample/$exit
      -- CP-element group 182: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(182)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(182)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(182) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_585_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_585_inst_ack_0, ack => maxPool4_CP_1841_elements(182)); -- 
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	319 
    -- CP-element group 183: 	384 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_update_completed_
      -- CP-element group 183: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_Update/ca
      -- CP-element group 183: 	 assign_stmt_417_to_assign_stmt_1457/slice_585_Update/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(183)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(183)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(183) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_585_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_585_inst_ack_1, ack => maxPool4_CP_1841_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	47 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_sample_start_
      -- CP-element group 184: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_Sample/rr
      -- CP-element group 184: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_Sample/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(184)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(184)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(184) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_589_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(184), ack => slice_589_inst_req_0); -- 
    maxPool4_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(186);
      gj_maxPool4_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: 	321 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_update_start_
      -- CP-element group 185: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_Update/$entry
      -- CP-element group 185: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(185)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(185)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(185) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_589_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(185), ack => slice_589_inst_req_1); -- 
    maxPool4_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(187) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	45 
    -- CP-element group 186: 	184 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_Sample/ra
      -- CP-element group 186: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_Sample/$exit
      -- CP-element group 186: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(186)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(186)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(186) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_589_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_589_inst_ack_0, ack => maxPool4_CP_1841_elements(186)); -- 
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	319 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	185 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_Update/$exit
      -- CP-element group 187: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_update_completed_
      -- CP-element group 187: 	 assign_stmt_417_to_assign_stmt_1457/slice_589_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(187)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(187)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(187) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_589_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_589_inst_ack_1, ack => maxPool4_CP_1841_elements(187)); -- 
    -- CP-element group 188:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	47 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	190 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_Sample/rr
      -- CP-element group 188: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_Sample/$entry
      -- CP-element group 188: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(188)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(188)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(188) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_593_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(188), ack => slice_593_inst_req_0); -- 
    maxPool4_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(190);
      gj_maxPool4_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: 	321 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_Update/cr
      -- CP-element group 189: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_Update/$entry
      -- CP-element group 189: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(189)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(189)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(189) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_593_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(189), ack => slice_593_inst_req_1); -- 
    maxPool4_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(191) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: marked-successors 
    -- CP-element group 190: 	45 
    -- CP-element group 190: 	188 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_Sample/ra
      -- CP-element group 190: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_Sample/$exit
      -- CP-element group 190: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(190)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(190)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(190) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_593_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_593_inst_ack_0, ack => maxPool4_CP_1841_elements(190)); -- 
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	319 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_Update/ca
      -- CP-element group 191: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_Update/$exit
      -- CP-element group 191: 	 assign_stmt_417_to_assign_stmt_1457/slice_593_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(191)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(191)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(191) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_593_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_593_inst_ack_1, ack => maxPool4_CP_1841_elements(191)); -- 
    -- CP-element group 192:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	47 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_Sample/$entry
      -- CP-element group 192: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_sample_start_
      -- CP-element group 192: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(192)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(192)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(192) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_597_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(192), ack => slice_597_inst_req_0); -- 
    maxPool4_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(194);
      gj_maxPool4_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: 	321 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_Update/$entry
      -- CP-element group 193: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_update_start_
      -- CP-element group 193: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(193)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(193)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(193) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_597_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(193), ack => slice_597_inst_req_1); -- 
    maxPool4_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(195) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	45 
    -- CP-element group 194: 	192 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_Sample/$exit
      -- CP-element group 194: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_sample_completed_
      -- CP-element group 194: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(194)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(194)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(194) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_597_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_597_inst_ack_0, ack => maxPool4_CP_1841_elements(194)); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	319 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_update_completed_
      -- CP-element group 195: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_Update/$exit
      -- CP-element group 195: 	 assign_stmt_417_to_assign_stmt_1457/slice_597_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(195)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(195)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(195) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_597_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_597_inst_ack_1, ack => maxPool4_CP_1841_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	47 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_Sample/rr
      -- CP-element group 196: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_Sample/$entry
      -- CP-element group 196: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(196)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(196)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(196) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_601_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(196), ack => slice_601_inst_req_0); -- 
    maxPool4_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(198);
      gj_maxPool4_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	199 
    -- CP-element group 197: 	340 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_Update/cr
      -- CP-element group 197: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_Update/$entry
      -- CP-element group 197: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(197)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(197)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(197) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_601_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(197), ack => slice_601_inst_req_1); -- 
    maxPool4_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(199) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	45 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_Sample/ra
      -- CP-element group 198: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_Sample/$exit
      -- CP-element group 198: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(198)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(198)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(198) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_601_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_601_inst_ack_0, ack => maxPool4_CP_1841_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	338 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	197 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_Update/$exit
      -- CP-element group 199: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_Update/ca
      -- CP-element group 199: 	 assign_stmt_417_to_assign_stmt_1457/slice_601_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(199)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(199)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(199) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_601_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_601_inst_ack_1, ack => maxPool4_CP_1841_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	47 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_Sample/rr
      -- CP-element group 200: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_Sample/$entry
      -- CP-element group 200: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(200)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(200)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(200) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_605_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(200), ack => slice_605_inst_req_0); -- 
    maxPool4_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(202);
      gj_maxPool4_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	203 
    -- CP-element group 201: 	340 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	203 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_Update/cr
      -- CP-element group 201: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_update_start_
      -- CP-element group 201: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_Update/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(201)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(201)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(201) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_605_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(201), ack => slice_605_inst_req_1); -- 
    maxPool4_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(203) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: successors 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	45 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_Sample/ra
      -- CP-element group 202: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_Sample/$exit
      -- CP-element group 202: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(202)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(202)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(202) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_605_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_605_inst_ack_0, ack => maxPool4_CP_1841_elements(202)); -- 
    -- CP-element group 203:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	201 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	338 
    -- CP-element group 203: marked-successors 
    -- CP-element group 203: 	201 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_Update/ca
      -- CP-element group 203: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_update_completed_
      -- CP-element group 203: 	 assign_stmt_417_to_assign_stmt_1457/slice_605_Update/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(203)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(203)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(203) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_605_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_605_inst_ack_1, ack => maxPool4_CP_1841_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	47 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	206 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_sample_start_
      -- CP-element group 204: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_Sample/rr
      -- CP-element group 204: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_Sample/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(204)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(204)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(204) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_609_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(204), ack => slice_609_inst_req_0); -- 
    maxPool4_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(206);
      gj_maxPool4_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: marked-predecessors 
    -- CP-element group 205: 	207 
    -- CP-element group 205: 	340 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_update_start_
      -- CP-element group 205: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_Update/$entry
      -- CP-element group 205: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(205)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(205)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(205) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_609_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(205), ack => slice_609_inst_req_1); -- 
    maxPool4_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(207) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	45 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_sample_completed_
      -- CP-element group 206: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_Sample/ra
      -- CP-element group 206: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_Sample/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(206)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(206)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(206) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_609_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_609_inst_ack_0, ack => maxPool4_CP_1841_elements(206)); -- 
    -- CP-element group 207:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	338 
    -- CP-element group 207: marked-successors 
    -- CP-element group 207: 	205 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_update_completed_
      -- CP-element group 207: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_Update/$exit
      -- CP-element group 207: 	 assign_stmt_417_to_assign_stmt_1457/slice_609_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(207)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(207)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(207) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_609_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_609_inst_ack_1, ack => maxPool4_CP_1841_elements(207)); -- 
    -- CP-element group 208:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	47 
    -- CP-element group 208: marked-predecessors 
    -- CP-element group 208: 	210 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_sample_start_
      -- CP-element group 208: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_Sample/rr
      -- CP-element group 208: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_Sample/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(208)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(208)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(208) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_613_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(208), ack => slice_613_inst_req_0); -- 
    maxPool4_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(210);
      gj_maxPool4_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: marked-predecessors 
    -- CP-element group 209: 	211 
    -- CP-element group 209: 	340 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_Update/$entry
      -- CP-element group 209: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_Update/cr
      -- CP-element group 209: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(209)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(209)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(209) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_613_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(209), ack => slice_613_inst_req_1); -- 
    maxPool4_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(211) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: marked-successors 
    -- CP-element group 210: 	45 
    -- CP-element group 210: 	208 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_sample_completed_
      -- CP-element group 210: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_Sample/ra
      -- CP-element group 210: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_Sample/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(210)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(210)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(210) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_613_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_613_inst_ack_0, ack => maxPool4_CP_1841_elements(210)); -- 
    -- CP-element group 211:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	338 
    -- CP-element group 211: marked-successors 
    -- CP-element group 211: 	209 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_Update/ca
      -- CP-element group 211: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_Update/$exit
      -- CP-element group 211: 	 assign_stmt_417_to_assign_stmt_1457/slice_613_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(211)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(211)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(211) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_613_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_613_inst_ack_1, ack => maxPool4_CP_1841_elements(211)); -- 
    -- CP-element group 212:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	47 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	214 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_Sample/rr
      -- CP-element group 212: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_sample_start_
      -- CP-element group 212: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_Sample/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(212)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(212)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(212) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_617_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(212), ack => slice_617_inst_req_0); -- 
    maxPool4_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(214);
      gj_maxPool4_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: marked-predecessors 
    -- CP-element group 213: 	215 
    -- CP-element group 213: 	359 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	215 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_update_start_
      -- CP-element group 213: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_Update/cr
      -- CP-element group 213: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_Update/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(213)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(213)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(213) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_617_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(213), ack => slice_617_inst_req_1); -- 
    maxPool4_cp_element_group_213: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_213"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(215) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_213 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(213), clk => clk, reset => reset); --
    end block;
    -- CP-element group 214:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214: marked-successors 
    -- CP-element group 214: 	45 
    -- CP-element group 214: 	212 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_Sample/ra
      -- CP-element group 214: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_sample_completed_
      -- CP-element group 214: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_Sample/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(214)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(214)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(214) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_617_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_617_inst_ack_0, ack => maxPool4_CP_1841_elements(214)); -- 
    -- CP-element group 215:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	213 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	357 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	213 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_update_completed_
      -- CP-element group 215: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_Update/ca
      -- CP-element group 215: 	 assign_stmt_417_to_assign_stmt_1457/slice_617_Update/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(215)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(215)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(215) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_617_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_617_inst_ack_1, ack => maxPool4_CP_1841_elements(215)); -- 
    -- CP-element group 216:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	47 
    -- CP-element group 216: marked-predecessors 
    -- CP-element group 216: 	218 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	218 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_Sample/$entry
      -- CP-element group 216: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_Sample/rr
      -- CP-element group 216: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(216)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(216)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(216) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_621_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(216), ack => slice_621_inst_req_0); -- 
    maxPool4_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(218);
      gj_maxPool4_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: 	359 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_Update/cr
      -- CP-element group 217: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_update_start_
      -- CP-element group 217: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_Update/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(217)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(217)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(217) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_621_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(217), ack => slice_621_inst_req_1); -- 
    maxPool4_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(219) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	45 
    -- CP-element group 218: 	216 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_Sample/$exit
      -- CP-element group 218: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_Sample/ra
      -- CP-element group 218: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(218)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(218)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(218) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_621_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_621_inst_ack_0, ack => maxPool4_CP_1841_elements(218)); -- 
    -- CP-element group 219:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	357 
    -- CP-element group 219: marked-successors 
    -- CP-element group 219: 	217 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_update_completed_
      -- CP-element group 219: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_Update/$exit
      -- CP-element group 219: 	 assign_stmt_417_to_assign_stmt_1457/slice_621_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(219)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(219)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(219) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_621_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_621_inst_ack_1, ack => maxPool4_CP_1841_elements(219)); -- 
    -- CP-element group 220:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	47 
    -- CP-element group 220: marked-predecessors 
    -- CP-element group 220: 	222 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_Sample/$entry
      -- CP-element group 220: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_sample_start_
      -- CP-element group 220: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(220)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(220)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(220) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_625_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(220), ack => slice_625_inst_req_0); -- 
    maxPool4_cp_element_group_220: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_220"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(222);
      gj_maxPool4_cp_element_group_220 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	223 
    -- CP-element group 221: 	359 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_update_start_
      -- CP-element group 221: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_Update/$entry
      -- CP-element group 221: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(221)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(221)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(221) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_625_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(221), ack => slice_625_inst_req_1); -- 
    maxPool4_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(223) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	45 
    -- CP-element group 222: 	220 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_sample_completed_
      -- CP-element group 222: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_Sample/$exit
      -- CP-element group 222: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(222)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(222)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(222) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_625_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_625_inst_ack_0, ack => maxPool4_CP_1841_elements(222)); -- 
    -- CP-element group 223:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	357 
    -- CP-element group 223: marked-successors 
    -- CP-element group 223: 	221 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_update_completed_
      -- CP-element group 223: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_Update/$exit
      -- CP-element group 223: 	 assign_stmt_417_to_assign_stmt_1457/slice_625_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(223)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(223)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(223) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_625_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_625_inst_ack_1, ack => maxPool4_CP_1841_elements(223)); -- 
    -- CP-element group 224:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	47 
    -- CP-element group 224: marked-predecessors 
    -- CP-element group 224: 	226 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	226 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_sample_start_
      -- CP-element group 224: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_Sample/$entry
      -- CP-element group 224: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(224)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(224)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(224) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_629_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(224), ack => slice_629_inst_req_0); -- 
    maxPool4_cp_element_group_224: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_224"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(226);
      gj_maxPool4_cp_element_group_224 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(224), clk => clk, reset => reset); --
    end block;
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	227 
    -- CP-element group 225: 	359 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_update_start_
      -- CP-element group 225: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_Update/$entry
      -- CP-element group 225: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(225)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(225)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(225) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_629_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(225), ack => slice_629_inst_req_1); -- 
    maxPool4_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(227) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	224 
    -- CP-element group 226: successors 
    -- CP-element group 226: marked-successors 
    -- CP-element group 226: 	45 
    -- CP-element group 226: 	224 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_sample_completed_
      -- CP-element group 226: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_Sample/$exit
      -- CP-element group 226: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(226)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(226)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(226) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_629_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_629_inst_ack_0, ack => maxPool4_CP_1841_elements(226)); -- 
    -- CP-element group 227:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	357 
    -- CP-element group 227: marked-successors 
    -- CP-element group 227: 	225 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_update_completed_
      -- CP-element group 227: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_Update/$exit
      -- CP-element group 227: 	 assign_stmt_417_to_assign_stmt_1457/slice_629_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(227)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(227)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(227) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_629_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_629_inst_ack_1, ack => maxPool4_CP_1841_elements(227)); -- 
    -- CP-element group 228:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	47 
    -- CP-element group 228: marked-predecessors 
    -- CP-element group 228: 	230 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_sample_start_
      -- CP-element group 228: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_Sample/$entry
      -- CP-element group 228: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(228)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(228)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(228) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_633_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(228), ack => slice_633_inst_req_0); -- 
    maxPool4_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(230);
      gj_maxPool4_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	231 
    -- CP-element group 229: 	378 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_update_start_
      -- CP-element group 229: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_Update/$entry
      -- CP-element group 229: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(229)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(229)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(229) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_633_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(229), ack => slice_633_inst_req_1); -- 
    maxPool4_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(231) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	45 
    -- CP-element group 230: 	228 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_sample_completed_
      -- CP-element group 230: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_Sample/$exit
      -- CP-element group 230: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(230)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(230)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(230) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_633_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_633_inst_ack_0, ack => maxPool4_CP_1841_elements(230)); -- 
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	376 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	229 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_update_completed_
      -- CP-element group 231: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_Update/$exit
      -- CP-element group 231: 	 assign_stmt_417_to_assign_stmt_1457/slice_633_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(231)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(231)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(231) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_633_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_633_inst_ack_1, ack => maxPool4_CP_1841_elements(231)); -- 
    -- CP-element group 232:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	47 
    -- CP-element group 232: marked-predecessors 
    -- CP-element group 232: 	234 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_sample_start_
      -- CP-element group 232: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_Sample/$entry
      -- CP-element group 232: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(232)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(232)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(232) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_637_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(232), ack => slice_637_inst_req_0); -- 
    maxPool4_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(234);
      gj_maxPool4_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: 	378 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_update_start_
      -- CP-element group 233: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_Update/$entry
      -- CP-element group 233: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(233)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(233)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(233) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_637_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(233), ack => slice_637_inst_req_1); -- 
    maxPool4_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(235) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: successors 
    -- CP-element group 234: marked-successors 
    -- CP-element group 234: 	45 
    -- CP-element group 234: 	232 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_sample_completed_
      -- CP-element group 234: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_Sample/$exit
      -- CP-element group 234: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(234)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(234)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(234) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_637_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_637_inst_ack_0, ack => maxPool4_CP_1841_elements(234)); -- 
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	376 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_update_completed_
      -- CP-element group 235: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_Update/$exit
      -- CP-element group 235: 	 assign_stmt_417_to_assign_stmt_1457/slice_637_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(235)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(235)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(235) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_637_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_637_inst_ack_1, ack => maxPool4_CP_1841_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	47 
    -- CP-element group 236: marked-predecessors 
    -- CP-element group 236: 	238 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	238 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_sample_start_
      -- CP-element group 236: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_Sample/$entry
      -- CP-element group 236: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(236)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(236)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(236) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_641_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(236), ack => slice_641_inst_req_0); -- 
    maxPool4_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(238);
      gj_maxPool4_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: 	378 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_update_start_
      -- CP-element group 237: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_Update/$entry
      -- CP-element group 237: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(237)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(237)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(237) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_641_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(237), ack => slice_641_inst_req_1); -- 
    maxPool4_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(239) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	236 
    -- CP-element group 238: successors 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	45 
    -- CP-element group 238: 	236 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_sample_completed_
      -- CP-element group 238: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_Sample/$exit
      -- CP-element group 238: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(238)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(238)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(238) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_641_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_641_inst_ack_0, ack => maxPool4_CP_1841_elements(238)); -- 
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	376 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_update_completed_
      -- CP-element group 239: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_Update/$exit
      -- CP-element group 239: 	 assign_stmt_417_to_assign_stmt_1457/slice_641_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(239)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(239)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(239) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_641_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_641_inst_ack_1, ack => maxPool4_CP_1841_elements(239)); -- 
    -- CP-element group 240:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	47 
    -- CP-element group 240: marked-predecessors 
    -- CP-element group 240: 	242 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_sample_start_
      -- CP-element group 240: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_Sample/$entry
      -- CP-element group 240: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(240)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(240)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(240) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_645_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(240), ack => slice_645_inst_req_0); -- 
    maxPool4_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(47) & maxPool4_CP_1841_elements(242);
      gj_maxPool4_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: 	378 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_update_start_
      -- CP-element group 241: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_Update/$entry
      -- CP-element group 241: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(241)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(241)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(241) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_645_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(241), ack => slice_645_inst_req_1); -- 
    maxPool4_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(243) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	240 
    -- CP-element group 242: successors 
    -- CP-element group 242: marked-successors 
    -- CP-element group 242: 	45 
    -- CP-element group 242: 	240 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_sample_completed_
      -- CP-element group 242: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_Sample/$exit
      -- CP-element group 242: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(242)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(242)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(242) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_645_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_645_inst_ack_0, ack => maxPool4_CP_1841_elements(242)); -- 
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	376 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_update_completed_
      -- CP-element group 243: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_Update/$exit
      -- CP-element group 243: 	 assign_stmt_417_to_assign_stmt_1457/slice_645_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(243)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(243)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(243) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_645_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_645_inst_ack_1, ack => maxPool4_CP_1841_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	51 
    -- CP-element group 244: marked-predecessors 
    -- CP-element group 244: 	246 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	246 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_sample_start_
      -- CP-element group 244: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_Sample/$entry
      -- CP-element group 244: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(244)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(244)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(244) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_649_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(244), ack => slice_649_inst_req_0); -- 
    maxPool4_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(246);
      gj_maxPool4_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: 	321 
    -- CP-element group 245: 	386 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_update_start_
      -- CP-element group 245: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_Update/$entry
      -- CP-element group 245: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(245)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(245)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(245) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_649_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(245), ack => slice_649_inst_req_1); -- 
    maxPool4_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(247) & maxPool4_CP_1841_elements(321) & maxPool4_CP_1841_elements(386);
      gj_maxPool4_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	244 
    -- CP-element group 246: successors 
    -- CP-element group 246: marked-successors 
    -- CP-element group 246: 	49 
    -- CP-element group 246: 	244 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_sample_completed_
      -- CP-element group 246: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_Sample/$exit
      -- CP-element group 246: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(246)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(246)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(246) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_649_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_649_inst_ack_0, ack => maxPool4_CP_1841_elements(246)); -- 
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	319 
    -- CP-element group 247: 	384 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_update_completed_
      -- CP-element group 247: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_Update/$exit
      -- CP-element group 247: 	 assign_stmt_417_to_assign_stmt_1457/slice_649_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(247)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(247)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(247) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_649_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_649_inst_ack_1, ack => maxPool4_CP_1841_elements(247)); -- 
    -- CP-element group 248:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	51 
    -- CP-element group 248: marked-predecessors 
    -- CP-element group 248: 	250 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_sample_start_
      -- CP-element group 248: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_Sample/$entry
      -- CP-element group 248: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(248)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(248)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(248) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_653_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(248), ack => slice_653_inst_req_0); -- 
    maxPool4_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(250);
      gj_maxPool4_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: 	321 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_update_start_
      -- CP-element group 249: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_Update/$entry
      -- CP-element group 249: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(249)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(249)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(249) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_653_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(249), ack => slice_653_inst_req_1); -- 
    maxPool4_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(251) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: marked-successors 
    -- CP-element group 250: 	49 
    -- CP-element group 250: 	248 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_sample_completed_
      -- CP-element group 250: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_Sample/$exit
      -- CP-element group 250: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(250)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(250)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(250) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_653_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_653_inst_ack_0, ack => maxPool4_CP_1841_elements(250)); -- 
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	319 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_update_completed_
      -- CP-element group 251: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_Update/$exit
      -- CP-element group 251: 	 assign_stmt_417_to_assign_stmt_1457/slice_653_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(251)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(251)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(251) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_653_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_653_inst_ack_1, ack => maxPool4_CP_1841_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	51 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_sample_start_
      -- CP-element group 252: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_Sample/$entry
      -- CP-element group 252: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(252)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(252)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(252) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_657_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(252), ack => slice_657_inst_req_0); -- 
    maxPool4_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(254);
      gj_maxPool4_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: 	321 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_update_start_
      -- CP-element group 253: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_Update/$entry
      -- CP-element group 253: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(253)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(253)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(253) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_657_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(253), ack => slice_657_inst_req_1); -- 
    maxPool4_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(255) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	49 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_sample_completed_
      -- CP-element group 254: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_Sample/$exit
      -- CP-element group 254: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(254)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(254)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(254) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_657_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_657_inst_ack_0, ack => maxPool4_CP_1841_elements(254)); -- 
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	319 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_update_completed_
      -- CP-element group 255: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_Update/$exit
      -- CP-element group 255: 	 assign_stmt_417_to_assign_stmt_1457/slice_657_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(255)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(255)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(255) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_657_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_657_inst_ack_1, ack => maxPool4_CP_1841_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	51 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_sample_start_
      -- CP-element group 256: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_Sample/$entry
      -- CP-element group 256: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(256)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(256)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(256) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_661_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(256), ack => slice_661_inst_req_0); -- 
    maxPool4_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(258);
      gj_maxPool4_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: 	321 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_update_start_
      -- CP-element group 257: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_Update/$entry
      -- CP-element group 257: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(257)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(257)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(257) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_661_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(257), ack => slice_661_inst_req_1); -- 
    maxPool4_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(259) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	49 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_sample_completed_
      -- CP-element group 258: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_Sample/$exit
      -- CP-element group 258: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(258)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(258)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(258) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_661_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_661_inst_ack_0, ack => maxPool4_CP_1841_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	319 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_update_completed_
      -- CP-element group 259: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_Update/$exit
      -- CP-element group 259: 	 assign_stmt_417_to_assign_stmt_1457/slice_661_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(259)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(259)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(259) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_661_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_661_inst_ack_1, ack => maxPool4_CP_1841_elements(259)); -- 
    -- CP-element group 260:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	51 
    -- CP-element group 260: marked-predecessors 
    -- CP-element group 260: 	262 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_sample_start_
      -- CP-element group 260: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_Sample/$entry
      -- CP-element group 260: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(260)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(260)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(260) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_665_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(260), ack => slice_665_inst_req_0); -- 
    maxPool4_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(262);
      gj_maxPool4_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: 	340 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_update_start_
      -- CP-element group 261: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_Update/$entry
      -- CP-element group 261: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(261)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(261)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(261) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_665_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(261), ack => slice_665_inst_req_1); -- 
    maxPool4_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(263) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262: marked-successors 
    -- CP-element group 262: 	49 
    -- CP-element group 262: 	260 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_sample_completed_
      -- CP-element group 262: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_Sample/$exit
      -- CP-element group 262: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(262)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(262)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(262) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_665_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_665_inst_ack_0, ack => maxPool4_CP_1841_elements(262)); -- 
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	338 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_update_completed_
      -- CP-element group 263: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_Update/$exit
      -- CP-element group 263: 	 assign_stmt_417_to_assign_stmt_1457/slice_665_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(263)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(263)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(263) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_665_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_665_inst_ack_1, ack => maxPool4_CP_1841_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	51 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	266 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_sample_start_
      -- CP-element group 264: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_Sample/$entry
      -- CP-element group 264: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(264)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(264)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(264) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_669_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(264), ack => slice_669_inst_req_0); -- 
    maxPool4_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(266);
      gj_maxPool4_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: 	340 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_update_start_
      -- CP-element group 265: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_Update/$entry
      -- CP-element group 265: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(265)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(265)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(265) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_669_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(265), ack => slice_669_inst_req_1); -- 
    maxPool4_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(267) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: marked-successors 
    -- CP-element group 266: 	49 
    -- CP-element group 266: 	264 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_sample_completed_
      -- CP-element group 266: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_Sample/$exit
      -- CP-element group 266: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(266)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(266)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(266) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_669_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_669_inst_ack_0, ack => maxPool4_CP_1841_elements(266)); -- 
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	338 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_update_completed_
      -- CP-element group 267: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_Update/$exit
      -- CP-element group 267: 	 assign_stmt_417_to_assign_stmt_1457/slice_669_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(267)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(267)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(267) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_669_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_669_inst_ack_1, ack => maxPool4_CP_1841_elements(267)); -- 
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	51 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	270 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_sample_start_
      -- CP-element group 268: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_Sample/$entry
      -- CP-element group 268: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(268)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(268)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(268) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_673_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(268), ack => slice_673_inst_req_0); -- 
    maxPool4_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(270);
      gj_maxPool4_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: 	340 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_update_start_
      -- CP-element group 269: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_Update/$entry
      -- CP-element group 269: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(269)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(269)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(269) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_673_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(269), ack => slice_673_inst_req_1); -- 
    maxPool4_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(271) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	49 
    -- CP-element group 270: 	268 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_sample_completed_
      -- CP-element group 270: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_Sample/$exit
      -- CP-element group 270: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(270)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(270)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(270) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_673_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_673_inst_ack_0, ack => maxPool4_CP_1841_elements(270)); -- 
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	338 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_update_completed_
      -- CP-element group 271: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_Update/$exit
      -- CP-element group 271: 	 assign_stmt_417_to_assign_stmt_1457/slice_673_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(271)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(271)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(271) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_673_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_673_inst_ack_1, ack => maxPool4_CP_1841_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	51 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_sample_start_
      -- CP-element group 272: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_Sample/$entry
      -- CP-element group 272: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(272)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(272)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(272) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_677_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(272), ack => slice_677_inst_req_0); -- 
    maxPool4_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(274);
      gj_maxPool4_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: 	340 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_update_start_
      -- CP-element group 273: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_Update/$entry
      -- CP-element group 273: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(273)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(273)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(273) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_677_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(273), ack => slice_677_inst_req_1); -- 
    maxPool4_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(275) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	49 
    -- CP-element group 274: 	272 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_sample_completed_
      -- CP-element group 274: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_Sample/$exit
      -- CP-element group 274: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(274)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(274)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(274) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_677_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_677_inst_ack_0, ack => maxPool4_CP_1841_elements(274)); -- 
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	338 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_update_completed_
      -- CP-element group 275: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_Update/$exit
      -- CP-element group 275: 	 assign_stmt_417_to_assign_stmt_1457/slice_677_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(275)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(275)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(275) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_677_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_677_inst_ack_1, ack => maxPool4_CP_1841_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	51 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_sample_start_
      -- CP-element group 276: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_Sample/$entry
      -- CP-element group 276: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(276)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(276)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(276) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_681_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(276), ack => slice_681_inst_req_0); -- 
    maxPool4_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(278);
      gj_maxPool4_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: 	359 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_update_start_
      -- CP-element group 277: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_Update/$entry
      -- CP-element group 277: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(277)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(277)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(277) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_681_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(277), ack => slice_681_inst_req_1); -- 
    maxPool4_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(279) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	49 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_sample_completed_
      -- CP-element group 278: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_Sample/$exit
      -- CP-element group 278: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(278)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(278)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(278) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_681_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_681_inst_ack_0, ack => maxPool4_CP_1841_elements(278)); -- 
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	357 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_update_completed_
      -- CP-element group 279: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_Update/$exit
      -- CP-element group 279: 	 assign_stmt_417_to_assign_stmt_1457/slice_681_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(279)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(279)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(279) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_681_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_681_inst_ack_1, ack => maxPool4_CP_1841_elements(279)); -- 
    -- CP-element group 280:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	51 
    -- CP-element group 280: marked-predecessors 
    -- CP-element group 280: 	282 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_sample_start_
      -- CP-element group 280: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_Sample/$entry
      -- CP-element group 280: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(280)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(280)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(280) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_685_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(280), ack => slice_685_inst_req_0); -- 
    maxPool4_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(282);
      gj_maxPool4_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	283 
    -- CP-element group 281: 	359 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_update_start_
      -- CP-element group 281: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_Update/$entry
      -- CP-element group 281: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(281)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(281)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(281) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_685_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(281), ack => slice_685_inst_req_1); -- 
    maxPool4_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(283) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: successors 
    -- CP-element group 282: marked-successors 
    -- CP-element group 282: 	49 
    -- CP-element group 282: 	280 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_sample_completed_
      -- CP-element group 282: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_Sample/$exit
      -- CP-element group 282: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(282)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(282)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(282) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_685_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_685_inst_ack_0, ack => maxPool4_CP_1841_elements(282)); -- 
    -- CP-element group 283:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	357 
    -- CP-element group 283: marked-successors 
    -- CP-element group 283: 	281 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_update_completed_
      -- CP-element group 283: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_Update/$exit
      -- CP-element group 283: 	 assign_stmt_417_to_assign_stmt_1457/slice_685_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(283)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(283)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(283) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_685_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_685_inst_ack_1, ack => maxPool4_CP_1841_elements(283)); -- 
    -- CP-element group 284:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	51 
    -- CP-element group 284: marked-predecessors 
    -- CP-element group 284: 	286 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	286 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_sample_start_
      -- CP-element group 284: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_Sample/$entry
      -- CP-element group 284: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(284)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(284)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(284) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_689_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(284), ack => slice_689_inst_req_0); -- 
    maxPool4_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(286);
      gj_maxPool4_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: 	359 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_update_start_
      -- CP-element group 285: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_Update/$entry
      -- CP-element group 285: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(285)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(285)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(285) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_689_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(285), ack => slice_689_inst_req_1); -- 
    maxPool4_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(287) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	284 
    -- CP-element group 286: successors 
    -- CP-element group 286: marked-successors 
    -- CP-element group 286: 	49 
    -- CP-element group 286: 	284 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_sample_completed_
      -- CP-element group 286: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_Sample/$exit
      -- CP-element group 286: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(286)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(286)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(286) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_689_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_689_inst_ack_0, ack => maxPool4_CP_1841_elements(286)); -- 
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	357 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	285 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_update_completed_
      -- CP-element group 287: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_Update/$exit
      -- CP-element group 287: 	 assign_stmt_417_to_assign_stmt_1457/slice_689_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(287)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(287)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(287) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_689_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_689_inst_ack_1, ack => maxPool4_CP_1841_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	51 
    -- CP-element group 288: marked-predecessors 
    -- CP-element group 288: 	290 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_sample_start_
      -- CP-element group 288: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_Sample/$entry
      -- CP-element group 288: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(288)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(288)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(288) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_693_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(288), ack => slice_693_inst_req_0); -- 
    maxPool4_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(290);
      gj_maxPool4_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: 	359 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_update_start_
      -- CP-element group 289: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_Update/$entry
      -- CP-element group 289: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(289)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(289)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(289) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_693_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(289), ack => slice_693_inst_req_1); -- 
    maxPool4_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(291) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: successors 
    -- CP-element group 290: marked-successors 
    -- CP-element group 290: 	49 
    -- CP-element group 290: 	288 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_sample_completed_
      -- CP-element group 290: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_Sample/$exit
      -- CP-element group 290: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(290)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(290)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(290) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_693_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_693_inst_ack_0, ack => maxPool4_CP_1841_elements(290)); -- 
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	357 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	289 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_update_completed_
      -- CP-element group 291: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_Update/$exit
      -- CP-element group 291: 	 assign_stmt_417_to_assign_stmt_1457/slice_693_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(291)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(291)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(291) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_693_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_693_inst_ack_1, ack => maxPool4_CP_1841_elements(291)); -- 
    -- CP-element group 292:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	51 
    -- CP-element group 292: marked-predecessors 
    -- CP-element group 292: 	294 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	294 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_sample_start_
      -- CP-element group 292: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_Sample/$entry
      -- CP-element group 292: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(292)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(292)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(292) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_697_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(292), ack => slice_697_inst_req_0); -- 
    maxPool4_cp_element_group_292: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_292"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(294);
      gj_maxPool4_cp_element_group_292 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(292), clk => clk, reset => reset); --
    end block;
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: 	378 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_update_start_
      -- CP-element group 293: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_Update/$entry
      -- CP-element group 293: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(293)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(293)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(293) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_697_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(293), ack => slice_697_inst_req_1); -- 
    maxPool4_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(295) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	292 
    -- CP-element group 294: successors 
    -- CP-element group 294: marked-successors 
    -- CP-element group 294: 	49 
    -- CP-element group 294: 	292 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_sample_completed_
      -- CP-element group 294: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_Sample/$exit
      -- CP-element group 294: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(294)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(294)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(294) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_697_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_697_inst_ack_0, ack => maxPool4_CP_1841_elements(294)); -- 
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	376 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_update_completed_
      -- CP-element group 295: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_Update/$exit
      -- CP-element group 295: 	 assign_stmt_417_to_assign_stmt_1457/slice_697_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(295)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(295)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(295) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_697_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_697_inst_ack_1, ack => maxPool4_CP_1841_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	51 
    -- CP-element group 296: marked-predecessors 
    -- CP-element group 296: 	298 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	298 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_sample_start_
      -- CP-element group 296: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_Sample/$entry
      -- CP-element group 296: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(296)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(296)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(296) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_701_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(296), ack => slice_701_inst_req_0); -- 
    maxPool4_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(298);
      gj_maxPool4_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: 	378 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_update_start_
      -- CP-element group 297: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_Update/$entry
      -- CP-element group 297: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(297)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(297)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(297) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_701_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(297), ack => slice_701_inst_req_1); -- 
    maxPool4_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(299) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	296 
    -- CP-element group 298: successors 
    -- CP-element group 298: marked-successors 
    -- CP-element group 298: 	49 
    -- CP-element group 298: 	296 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_sample_completed_
      -- CP-element group 298: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_Sample/$exit
      -- CP-element group 298: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(298)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(298)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(298) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_701_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_701_inst_ack_0, ack => maxPool4_CP_1841_elements(298)); -- 
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	376 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_update_completed_
      -- CP-element group 299: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_Update/$exit
      -- CP-element group 299: 	 assign_stmt_417_to_assign_stmt_1457/slice_701_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(299)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(299)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(299) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_701_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_701_inst_ack_1, ack => maxPool4_CP_1841_elements(299)); -- 
    -- CP-element group 300:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	51 
    -- CP-element group 300: marked-predecessors 
    -- CP-element group 300: 	302 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	302 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_sample_start_
      -- CP-element group 300: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_Sample/$entry
      -- CP-element group 300: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(300)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(300)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(300) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_705_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(300), ack => slice_705_inst_req_0); -- 
    maxPool4_cp_element_group_300: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_300"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(302);
      gj_maxPool4_cp_element_group_300 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(300), clk => clk, reset => reset); --
    end block;
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: 	378 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_Update/$entry
      -- CP-element group 301: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_Update/cr
      -- CP-element group 301: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(301)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(301)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(301) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_705_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(301), ack => slice_705_inst_req_1); -- 
    maxPool4_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(303) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	300 
    -- CP-element group 302: successors 
    -- CP-element group 302: marked-successors 
    -- CP-element group 302: 	49 
    -- CP-element group 302: 	300 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_sample_completed_
      -- CP-element group 302: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_Sample/$exit
      -- CP-element group 302: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(302)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(302)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(302) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_705_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_705_inst_ack_0, ack => maxPool4_CP_1841_elements(302)); -- 
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	376 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	301 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_Update/$exit
      -- CP-element group 303: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_Update/ca
      -- CP-element group 303: 	 assign_stmt_417_to_assign_stmt_1457/slice_705_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(303)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(303)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(303) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_705_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_705_inst_ack_1, ack => maxPool4_CP_1841_elements(303)); -- 
    -- CP-element group 304:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	51 
    -- CP-element group 304: marked-predecessors 
    -- CP-element group 304: 	306 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	306 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_sample_start_
      -- CP-element group 304: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_Sample/$entry
      -- CP-element group 304: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(304)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(304)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(304) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_709_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(304), ack => slice_709_inst_req_0); -- 
    maxPool4_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(51) & maxPool4_CP_1841_elements(306);
      gj_maxPool4_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: 	378 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_update_start_
      -- CP-element group 305: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_Update/$entry
      -- CP-element group 305: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(305)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(305)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(305) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_709_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(305), ack => slice_709_inst_req_1); -- 
    maxPool4_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(307) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	304 
    -- CP-element group 306: successors 
    -- CP-element group 306: marked-successors 
    -- CP-element group 306: 	49 
    -- CP-element group 306: 	304 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_sample_completed_
      -- CP-element group 306: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_Sample/$exit
      -- CP-element group 306: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(306)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(306)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(306) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_709_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_709_inst_ack_0, ack => maxPool4_CP_1841_elements(306)); -- 
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	376 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_update_completed_
      -- CP-element group 307: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_Update/$exit
      -- CP-element group 307: 	 assign_stmt_417_to_assign_stmt_1457/slice_709_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(307)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(307)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(307) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:slice_709_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_709_inst_ack_1, ack => maxPool4_CP_1841_elements(307)); -- 
    -- CP-element group 308:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	312 
    -- CP-element group 308: marked-predecessors 
    -- CP-element group 308: 	313 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	313 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_sample_start_
      -- CP-element group 308: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_request/$entry
      -- CP-element group 308: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_request/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(308)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(308)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(308) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1357_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(308), ack => addr_of_1357_final_reg_req_0); -- 
    maxPool4_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(312) & maxPool4_CP_1841_elements(313);
      gj_maxPool4_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	1 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	314 
    -- CP-element group 309: 	317 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	314 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_update_start_
      -- CP-element group 309: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_complete/$entry
      -- CP-element group 309: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_complete/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(309)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(309)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(309) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1357_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(309), ack => addr_of_1357_final_reg_req_1); -- 
    maxPool4_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(314) & maxPool4_CP_1841_elements(317);
      gj_maxPool4_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	1 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: 	313 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_final_index_sum_regn_update_start
      -- CP-element group 310: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_final_index_sum_regn_Update/$entry
      -- CP-element group 310: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_final_index_sum_regn_Update/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(310)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(310)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(310) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1356_index_offset_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(310), ack => array_obj_ref_1356_index_offset_req_1); -- 
    maxPool4_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(312) & maxPool4_CP_1841_elements(313);
      gj_maxPool4_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	1 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	391 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	2 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_final_index_sum_regn_sample_complete
      -- CP-element group 311: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_final_index_sum_regn_Sample/$exit
      -- CP-element group 311: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(311)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(311)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(311) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1356_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1356_index_offset_ack_0, ack => maxPool4_CP_1841_elements(311)); -- 
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	308 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	310 
    -- CP-element group 312:  members (8) 
      -- CP-element group 312: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_root_address_calculated
      -- CP-element group 312: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_offset_calculated
      -- CP-element group 312: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_final_index_sum_regn_Update/$exit
      -- CP-element group 312: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_final_index_sum_regn_Update/ack
      -- CP-element group 312: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_base_plus_offset/$entry
      -- CP-element group 312: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_base_plus_offset/$exit
      -- CP-element group 312: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_base_plus_offset/sum_rename_req
      -- CP-element group 312: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1356_base_plus_offset/sum_rename_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(312)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(312)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(312) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1356_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1356_index_offset_ack_1, ack => maxPool4_CP_1841_elements(312)); -- 
    -- CP-element group 313:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	308 
    -- CP-element group 313: successors 
    -- CP-element group 313: marked-successors 
    -- CP-element group 313: 	308 
    -- CP-element group 313: 	310 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_sample_completed_
      -- CP-element group 313: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_request/$exit
      -- CP-element group 313: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_request/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(313)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(313)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(313) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1357_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1357_final_reg_ack_0, ack => maxPool4_CP_1841_elements(313)); -- 
    -- CP-element group 314:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	309 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314: marked-successors 
    -- CP-element group 314: 	309 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_update_completed_
      -- CP-element group 314: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_complete/$exit
      -- CP-element group 314: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1357_complete/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(314)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(314)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(314) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1357_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1357_final_reg_ack_1, ack => maxPool4_CP_1841_elements(314)); -- 
    -- CP-element group 315:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: marked-predecessors 
    -- CP-element group 315: 	317 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_sample_start_
      -- CP-element group 315: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_Sample/$entry
      -- CP-element group 315: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_Sample/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(315)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(315)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(315) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr5_1359_delayed_8_0_1359_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(315), ack => W_myptr5_1359_delayed_8_0_1359_inst_req_0); -- 
    maxPool4_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(314) & maxPool4_CP_1841_elements(317);
      gj_maxPool4_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: marked-predecessors 
    -- CP-element group 316: 	318 
    -- CP-element group 316: 	325 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	318 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_update_start_
      -- CP-element group 316: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_Update/$entry
      -- CP-element group 316: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_Update/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(316)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(316)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(316) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr5_1359_delayed_8_0_1359_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(316), ack => W_myptr5_1359_delayed_8_0_1359_inst_req_1); -- 
    maxPool4_cp_element_group_316: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_316"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(318) & maxPool4_CP_1841_elements(325);
      gj_maxPool4_cp_element_group_316 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(316), clk => clk, reset => reset); --
    end block;
    -- CP-element group 317:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: successors 
    -- CP-element group 317: marked-successors 
    -- CP-element group 317: 	309 
    -- CP-element group 317: 	315 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_sample_completed_
      -- CP-element group 317: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_Sample/$exit
      -- CP-element group 317: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_Sample/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(317)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(317)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(317) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr5_1359_delayed_8_0_1359_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr5_1359_delayed_8_0_1359_inst_ack_0, ack => maxPool4_CP_1841_elements(317)); -- 
    -- CP-element group 318:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	316 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	323 
    -- CP-element group 318: marked-successors 
    -- CP-element group 318: 	316 
    -- CP-element group 318:  members (19) 
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_word_addrgen/root_register_ack
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_word_addrgen/root_register_req
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_word_addrgen/$exit
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_word_addrgen/$entry
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_update_completed_
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_Update/$exit
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1361_Update/ack
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_base_address_calculated
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_word_address_calculated
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_root_address_calculated
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_base_address_resized
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_base_addr_resize/$entry
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_base_addr_resize/$exit
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_base_addr_resize/base_resize_req
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_base_addr_resize/base_resize_ack
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_base_plus_offset/$entry
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_base_plus_offset/$exit
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_base_plus_offset/sum_rename_req
      -- CP-element group 318: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_base_plus_offset/sum_rename_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(318)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(318)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(318) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr5_1359_delayed_8_0_1359_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr5_1359_delayed_8_0_1359_inst_ack_1, ack => maxPool4_CP_1841_elements(318)); -- 
    -- CP-element group 319:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	55 
    -- CP-element group 319: 	59 
    -- CP-element group 319: 	63 
    -- CP-element group 319: 	67 
    -- CP-element group 319: 	119 
    -- CP-element group 319: 	123 
    -- CP-element group 319: 	127 
    -- CP-element group 319: 	131 
    -- CP-element group 319: 	183 
    -- CP-element group 319: 	187 
    -- CP-element group 319: 	191 
    -- CP-element group 319: 	195 
    -- CP-element group 319: 	247 
    -- CP-element group 319: 	251 
    -- CP-element group 319: 	255 
    -- CP-element group 319: 	259 
    -- CP-element group 319: marked-predecessors 
    -- CP-element group 319: 	321 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_sample_start_
      -- CP-element group 319: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_Sample/$entry
      -- CP-element group 319: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(319)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(319)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(319) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1374_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(319), ack => CONCAT_u32_u64_1374_inst_req_0); -- 
    maxPool4_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(55) & maxPool4_CP_1841_elements(59) & maxPool4_CP_1841_elements(63) & maxPool4_CP_1841_elements(67) & maxPool4_CP_1841_elements(119) & maxPool4_CP_1841_elements(123) & maxPool4_CP_1841_elements(127) & maxPool4_CP_1841_elements(131) & maxPool4_CP_1841_elements(183) & maxPool4_CP_1841_elements(187) & maxPool4_CP_1841_elements(191) & maxPool4_CP_1841_elements(195) & maxPool4_CP_1841_elements(247) & maxPool4_CP_1841_elements(251) & maxPool4_CP_1841_elements(255) & maxPool4_CP_1841_elements(259) & maxPool4_CP_1841_elements(321);
      gj_maxPool4_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: marked-predecessors 
    -- CP-element group 320: 	322 
    -- CP-element group 320: 	325 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	322 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_update_start_
      -- CP-element group 320: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_Update/$entry
      -- CP-element group 320: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(320)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(320)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(320) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1374_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(320), ack => CONCAT_u32_u64_1374_inst_req_1); -- 
    maxPool4_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(322) & maxPool4_CP_1841_elements(325);
      gj_maxPool4_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321: marked-successors 
    -- CP-element group 321: 	53 
    -- CP-element group 321: 	57 
    -- CP-element group 321: 	61 
    -- CP-element group 321: 	65 
    -- CP-element group 321: 	117 
    -- CP-element group 321: 	121 
    -- CP-element group 321: 	125 
    -- CP-element group 321: 	129 
    -- CP-element group 321: 	181 
    -- CP-element group 321: 	185 
    -- CP-element group 321: 	189 
    -- CP-element group 321: 	193 
    -- CP-element group 321: 	245 
    -- CP-element group 321: 	249 
    -- CP-element group 321: 	253 
    -- CP-element group 321: 	257 
    -- CP-element group 321: 	319 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_sample_completed_
      -- CP-element group 321: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_Sample/$exit
      -- CP-element group 321: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(321)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(321)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(321) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1374_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1374_inst_ack_0, ack => maxPool4_CP_1841_elements(321)); -- 
    -- CP-element group 322:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	320 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322: marked-successors 
    -- CP-element group 322: 	320 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_update_completed_
      -- CP-element group 322: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_Update/$exit
      -- CP-element group 322: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1374_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(322)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(322)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(322) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1374_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1374_inst_ack_1, ack => maxPool4_CP_1841_elements(322)); -- 
    -- CP-element group 323:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	318 
    -- CP-element group 323: 	322 
    -- CP-element group 323: marked-predecessors 
    -- CP-element group 323: 	325 
    -- CP-element group 323: 	382 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (9) 
      -- CP-element group 323: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/word_access_start/word_0/rr
      -- CP-element group 323: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/word_access_start/word_0/$entry
      -- CP-element group 323: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/word_access_start/$entry
      -- CP-element group 323: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/ptr_deref_1363_Split/split_ack
      -- CP-element group 323: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/ptr_deref_1363_Split/split_req
      -- CP-element group 323: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/ptr_deref_1363_Split/$exit
      -- CP-element group 323: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/ptr_deref_1363_Split/$entry
      -- CP-element group 323: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/$entry
      -- CP-element group 323: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(323)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(323)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(323) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1363_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(323), ack => ptr_deref_1363_store_0_req_0); -- 
    maxPool4_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(318) & maxPool4_CP_1841_elements(322) & maxPool4_CP_1841_elements(325) & maxPool4_CP_1841_elements(382);
      gj_maxPool4_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: marked-predecessors 
    -- CP-element group 324: 	326 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (5) 
      -- CP-element group 324: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Update/word_access_complete/word_0/cr
      -- CP-element group 324: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Update/word_access_complete/word_0/$entry
      -- CP-element group 324: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Update/word_access_complete/$entry
      -- CP-element group 324: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Update/$entry
      -- CP-element group 324: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(324)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(324)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(324) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1363_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(324), ack => ptr_deref_1363_store_0_req_1); -- 
    maxPool4_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_1841_elements(326);
      gj_maxPool4_cp_element_group_324 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	388 
    -- CP-element group 325: marked-successors 
    -- CP-element group 325: 	316 
    -- CP-element group 325: 	320 
    -- CP-element group 325: 	323 
    -- CP-element group 325:  members (5) 
      -- CP-element group 325: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/word_access_start/word_0/ra
      -- CP-element group 325: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/word_access_start/word_0/$exit
      -- CP-element group 325: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/word_access_start/$exit
      -- CP-element group 325: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Sample/$exit
      -- CP-element group 325: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(325)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(325)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(325) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1363_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1363_store_0_ack_0, ack => maxPool4_CP_1841_elements(325)); -- 
    -- CP-element group 326:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	391 
    -- CP-element group 326: marked-successors 
    -- CP-element group 326: 	324 
    -- CP-element group 326:  members (5) 
      -- CP-element group 326: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Update/word_access_complete/word_0/ca
      -- CP-element group 326: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Update/word_access_complete/word_0/$exit
      -- CP-element group 326: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Update/word_access_complete/$exit
      -- CP-element group 326: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_Update/$exit
      -- CP-element group 326: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(326)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(326)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(326) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1363_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1363_store_0_ack_1, ack => maxPool4_CP_1841_elements(326)); -- 
    -- CP-element group 327:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	331 
    -- CP-element group 327: marked-predecessors 
    -- CP-element group 327: 	332 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	332 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_sample_start_
      -- CP-element group 327: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_request/req
      -- CP-element group 327: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_request/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(327)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(327)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(327) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1383_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(327), ack => addr_of_1383_final_reg_req_0); -- 
    maxPool4_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(331) & maxPool4_CP_1841_elements(332);
      gj_maxPool4_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	1 
    -- CP-element group 328: marked-predecessors 
    -- CP-element group 328: 	333 
    -- CP-element group 328: 	336 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	333 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_update_start_
      -- CP-element group 328: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_complete/req
      -- CP-element group 328: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_complete/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(328)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(328)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(328) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1383_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(328), ack => addr_of_1383_final_reg_req_1); -- 
    maxPool4_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(333) & maxPool4_CP_1841_elements(336);
      gj_maxPool4_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	1 
    -- CP-element group 329: marked-predecessors 
    -- CP-element group 329: 	331 
    -- CP-element group 329: 	332 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_final_index_sum_regn_update_start
      -- CP-element group 329: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_final_index_sum_regn_Update/req
      -- CP-element group 329: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_final_index_sum_regn_Update/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(329)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(329)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(329) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1382_index_offset_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(329), ack => array_obj_ref_1382_index_offset_req_1); -- 
    maxPool4_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(331) & maxPool4_CP_1841_elements(332);
      gj_maxPool4_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	1 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	391 
    -- CP-element group 330: marked-successors 
    -- CP-element group 330: 	2 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_final_index_sum_regn_sample_complete
      -- CP-element group 330: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_final_index_sum_regn_Sample/ack
      -- CP-element group 330: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_final_index_sum_regn_Sample/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(330)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(330)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(330) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1382_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1382_index_offset_ack_0, ack => maxPool4_CP_1841_elements(330)); -- 
    -- CP-element group 331:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	327 
    -- CP-element group 331: marked-successors 
    -- CP-element group 331: 	329 
    -- CP-element group 331:  members (8) 
      -- CP-element group 331: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_root_address_calculated
      -- CP-element group 331: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_offset_calculated
      -- CP-element group 331: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_base_plus_offset/sum_rename_ack
      -- CP-element group 331: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_base_plus_offset/sum_rename_req
      -- CP-element group 331: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_base_plus_offset/$exit
      -- CP-element group 331: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_base_plus_offset/$entry
      -- CP-element group 331: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_final_index_sum_regn_Update/ack
      -- CP-element group 331: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1382_final_index_sum_regn_Update/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(331)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(331)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(331) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1382_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1382_index_offset_ack_1, ack => maxPool4_CP_1841_elements(331)); -- 
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	327 
    -- CP-element group 332: successors 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	327 
    -- CP-element group 332: 	329 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_sample_completed_
      -- CP-element group 332: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_request/ack
      -- CP-element group 332: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_request/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(332)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(332)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(332) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1383_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1383_final_reg_ack_0, ack => maxPool4_CP_1841_elements(332)); -- 
    -- CP-element group 333:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	328 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333: marked-successors 
    -- CP-element group 333: 	328 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_update_completed_
      -- CP-element group 333: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_complete/ack
      -- CP-element group 333: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1383_complete/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(333)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(333)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(333) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1383_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1383_final_reg_ack_1, ack => maxPool4_CP_1841_elements(333)); -- 
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_Sample/req
      -- CP-element group 334: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_Sample/$entry
      -- CP-element group 334: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(334)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(334)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(334) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr6_1382_delayed_8_0_1385_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(334), ack => W_myptr6_1382_delayed_8_0_1385_inst_req_0); -- 
    maxPool4_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(333) & maxPool4_CP_1841_elements(336);
      gj_maxPool4_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: marked-predecessors 
    -- CP-element group 335: 	337 
    -- CP-element group 335: 	344 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_Update/$entry
      -- CP-element group 335: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_Update/req
      -- CP-element group 335: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(335)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(335)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(335) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr6_1382_delayed_8_0_1385_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(335), ack => W_myptr6_1382_delayed_8_0_1385_inst_req_1); -- 
    maxPool4_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(337) & maxPool4_CP_1841_elements(344);
      gj_maxPool4_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	328 
    -- CP-element group 336: 	334 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_Sample/ack
      -- CP-element group 336: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_Sample/$exit
      -- CP-element group 336: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(336)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(336)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(336) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr6_1382_delayed_8_0_1385_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr6_1382_delayed_8_0_1385_inst_ack_0, ack => maxPool4_CP_1841_elements(336)); -- 
    -- CP-element group 337:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	342 
    -- CP-element group 337: marked-successors 
    -- CP-element group 337: 	335 
    -- CP-element group 337:  members (19) 
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_base_address_calculated
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_Update/$exit
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_Update/ack
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_base_plus_offset/$exit
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_base_plus_offset/sum_rename_req
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_base_plus_offset/sum_rename_ack
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_word_address_calculated
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_root_address_calculated
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_base_address_resized
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_base_addr_resize/$entry
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_word_addrgen/$entry
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_base_addr_resize/$exit
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_base_addr_resize/base_resize_req
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_word_addrgen/$exit
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_base_addr_resize/base_resize_ack
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_base_plus_offset/$entry
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1387_update_completed_
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_word_addrgen/root_register_ack
      -- CP-element group 337: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_word_addrgen/root_register_req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(337)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(337)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(337) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr6_1382_delayed_8_0_1385_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr6_1382_delayed_8_0_1385_inst_ack_1, ack => maxPool4_CP_1841_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	71 
    -- CP-element group 338: 	75 
    -- CP-element group 338: 	79 
    -- CP-element group 338: 	83 
    -- CP-element group 338: 	135 
    -- CP-element group 338: 	139 
    -- CP-element group 338: 	143 
    -- CP-element group 338: 	147 
    -- CP-element group 338: 	199 
    -- CP-element group 338: 	203 
    -- CP-element group 338: 	207 
    -- CP-element group 338: 	211 
    -- CP-element group 338: 	263 
    -- CP-element group 338: 	267 
    -- CP-element group 338: 	271 
    -- CP-element group 338: 	275 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_sample_start_
      -- CP-element group 338: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_Sample/$entry
      -- CP-element group 338: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(338)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(338)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(338) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1400_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(338), ack => CONCAT_u32_u64_1400_inst_req_0); -- 
    maxPool4_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(71) & maxPool4_CP_1841_elements(75) & maxPool4_CP_1841_elements(79) & maxPool4_CP_1841_elements(83) & maxPool4_CP_1841_elements(135) & maxPool4_CP_1841_elements(139) & maxPool4_CP_1841_elements(143) & maxPool4_CP_1841_elements(147) & maxPool4_CP_1841_elements(199) & maxPool4_CP_1841_elements(203) & maxPool4_CP_1841_elements(207) & maxPool4_CP_1841_elements(211) & maxPool4_CP_1841_elements(263) & maxPool4_CP_1841_elements(267) & maxPool4_CP_1841_elements(271) & maxPool4_CP_1841_elements(275) & maxPool4_CP_1841_elements(340);
      gj_maxPool4_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	341 
    -- CP-element group 339: 	344 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_update_start_
      -- CP-element group 339: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_Update/$entry
      -- CP-element group 339: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(339)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(339)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(339) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1400_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(339), ack => CONCAT_u32_u64_1400_inst_req_1); -- 
    maxPool4_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(341) & maxPool4_CP_1841_elements(344);
      gj_maxPool4_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	69 
    -- CP-element group 340: 	73 
    -- CP-element group 340: 	77 
    -- CP-element group 340: 	81 
    -- CP-element group 340: 	133 
    -- CP-element group 340: 	137 
    -- CP-element group 340: 	141 
    -- CP-element group 340: 	145 
    -- CP-element group 340: 	197 
    -- CP-element group 340: 	201 
    -- CP-element group 340: 	205 
    -- CP-element group 340: 	209 
    -- CP-element group 340: 	261 
    -- CP-element group 340: 	265 
    -- CP-element group 340: 	269 
    -- CP-element group 340: 	273 
    -- CP-element group 340: 	338 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_sample_completed_
      -- CP-element group 340: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_Sample/$exit
      -- CP-element group 340: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(340)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(340)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(340) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1400_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1400_inst_ack_0, ack => maxPool4_CP_1841_elements(340)); -- 
    -- CP-element group 341:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341: marked-successors 
    -- CP-element group 341: 	339 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_update_completed_
      -- CP-element group 341: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_Update/$exit
      -- CP-element group 341: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1400_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(341)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(341)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(341) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1400_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1400_inst_ack_1, ack => maxPool4_CP_1841_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	337 
    -- CP-element group 342: 	341 
    -- CP-element group 342: 	388 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (9) 
      -- CP-element group 342: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_sample_start_
      -- CP-element group 342: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/word_access_start/word_0/rr
      -- CP-element group 342: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/word_access_start/word_0/$entry
      -- CP-element group 342: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/word_access_start/$entry
      -- CP-element group 342: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/ptr_deref_1389_Split/split_ack
      -- CP-element group 342: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/ptr_deref_1389_Split/split_req
      -- CP-element group 342: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/ptr_deref_1389_Split/$exit
      -- CP-element group 342: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/ptr_deref_1389_Split/$entry
      -- CP-element group 342: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(342)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(342)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(342) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1389_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(342), ack => ptr_deref_1389_store_0_req_0); -- 
    maxPool4_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(337) & maxPool4_CP_1841_elements(341) & maxPool4_CP_1841_elements(388) & maxPool4_CP_1841_elements(344);
      gj_maxPool4_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	345 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343:  members (5) 
      -- CP-element group 343: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Update/word_access_complete/word_0/cr
      -- CP-element group 343: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Update/word_access_complete/word_0/$entry
      -- CP-element group 343: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Update/word_access_complete/$entry
      -- CP-element group 343: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Update/$entry
      -- CP-element group 343: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(343)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(343)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(343) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1389_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(343), ack => ptr_deref_1389_store_0_req_1); -- 
    maxPool4_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_1841_elements(345);
      gj_maxPool4_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	389 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	335 
    -- CP-element group 344: 	339 
    -- CP-element group 344: 	342 
    -- CP-element group 344:  members (5) 
      -- CP-element group 344: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_sample_completed_
      -- CP-element group 344: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/word_access_start/word_0/ra
      -- CP-element group 344: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/word_access_start/word_0/$exit
      -- CP-element group 344: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/word_access_start/$exit
      -- CP-element group 344: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Sample/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(344)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(344)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(344) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1389_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1389_store_0_ack_0, ack => maxPool4_CP_1841_elements(344)); -- 
    -- CP-element group 345:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	391 
    -- CP-element group 345: marked-successors 
    -- CP-element group 345: 	343 
    -- CP-element group 345:  members (5) 
      -- CP-element group 345: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_update_completed_
      -- CP-element group 345: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Update/word_access_complete/word_0/ca
      -- CP-element group 345: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Update/word_access_complete/word_0/$exit
      -- CP-element group 345: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Update/word_access_complete/$exit
      -- CP-element group 345: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_Update/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(345)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(345)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(345) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1389_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1389_store_0_ack_1, ack => maxPool4_CP_1841_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	350 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	351 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	351 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_sample_start_
      -- CP-element group 346: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_request/req
      -- CP-element group 346: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_request/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(346)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(346)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(346) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1409_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(346), ack => addr_of_1409_final_reg_req_0); -- 
    maxPool4_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(350) & maxPool4_CP_1841_elements(351);
      gj_maxPool4_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	1 
    -- CP-element group 347: marked-predecessors 
    -- CP-element group 347: 	352 
    -- CP-element group 347: 	355 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	352 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_complete/req
      -- CP-element group 347: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_update_start_
      -- CP-element group 347: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_complete/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(347)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(347)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(347) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1409_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(347), ack => addr_of_1409_final_reg_req_1); -- 
    maxPool4_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(352) & maxPool4_CP_1841_elements(355);
      gj_maxPool4_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	1 
    -- CP-element group 348: marked-predecessors 
    -- CP-element group 348: 	350 
    -- CP-element group 348: 	351 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	350 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_final_index_sum_regn_Update/req
      -- CP-element group 348: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_final_index_sum_regn_Update/$entry
      -- CP-element group 348: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_final_index_sum_regn_update_start
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(348)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(348)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(348) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1408_index_offset_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(348), ack => array_obj_ref_1408_index_offset_req_1); -- 
    maxPool4_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(350) & maxPool4_CP_1841_elements(351);
      gj_maxPool4_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	1 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	391 
    -- CP-element group 349: marked-successors 
    -- CP-element group 349: 	2 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_final_index_sum_regn_Sample/ack
      -- CP-element group 349: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_final_index_sum_regn_Sample/$exit
      -- CP-element group 349: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_final_index_sum_regn_sample_complete
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(349)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(349)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(349) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1408_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1408_index_offset_ack_0, ack => maxPool4_CP_1841_elements(349)); -- 
    -- CP-element group 350:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	348 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	346 
    -- CP-element group 350: marked-successors 
    -- CP-element group 350: 	348 
    -- CP-element group 350:  members (8) 
      -- CP-element group 350: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_final_index_sum_regn_Update/ack
      -- CP-element group 350: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_base_plus_offset/$entry
      -- CP-element group 350: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_base_plus_offset/$exit
      -- CP-element group 350: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_base_plus_offset/sum_rename_req
      -- CP-element group 350: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_final_index_sum_regn_Update/$exit
      -- CP-element group 350: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_offset_calculated
      -- CP-element group 350: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_root_address_calculated
      -- CP-element group 350: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1408_base_plus_offset/sum_rename_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(350)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(350)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(350) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1408_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1408_index_offset_ack_1, ack => maxPool4_CP_1841_elements(350)); -- 
    -- CP-element group 351:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	346 
    -- CP-element group 351: successors 
    -- CP-element group 351: marked-successors 
    -- CP-element group 351: 	346 
    -- CP-element group 351: 	348 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_sample_completed_
      -- CP-element group 351: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_request/ack
      -- CP-element group 351: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_request/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(351)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(351)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(351) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1409_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1409_final_reg_ack_0, ack => maxPool4_CP_1841_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	347 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	347 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_complete/ack
      -- CP-element group 352: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_update_completed_
      -- CP-element group 352: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1409_complete/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(352)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(352)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(352) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1409_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1409_final_reg_ack_1, ack => maxPool4_CP_1841_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: marked-predecessors 
    -- CP-element group 353: 	355 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_sample_start_
      -- CP-element group 353: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_Sample/$entry
      -- CP-element group 353: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_Sample/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(353)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(353)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(353) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr7_1405_delayed_8_0_1411_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(353), ack => W_myptr7_1405_delayed_8_0_1411_inst_req_0); -- 
    maxPool4_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(352) & maxPool4_CP_1841_elements(355);
      gj_maxPool4_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: 	363 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_update_start_
      -- CP-element group 354: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_Update/req
      -- CP-element group 354: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_Update/$entry
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(354)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(354)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(354) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr7_1405_delayed_8_0_1411_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(354), ack => W_myptr7_1405_delayed_8_0_1411_inst_req_1); -- 
    maxPool4_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(356) & maxPool4_CP_1841_elements(363);
      gj_maxPool4_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355: marked-successors 
    -- CP-element group 355: 	347 
    -- CP-element group 355: 	353 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_sample_completed_
      -- CP-element group 355: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_Sample/$exit
      -- CP-element group 355: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_Sample/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(355)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(355)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(355) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr7_1405_delayed_8_0_1411_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr7_1405_delayed_8_0_1411_inst_ack_0, ack => maxPool4_CP_1841_elements(355)); -- 
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	361 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (19) 
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_base_address_calculated
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_word_address_calculated
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_root_address_calculated
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_base_address_resized
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_base_addr_resize/$entry
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_word_addrgen/$exit
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_base_addr_resize/$exit
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_base_addr_resize/base_resize_req
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_base_addr_resize/base_resize_ack
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_base_plus_offset/$entry
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_update_completed_
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_base_plus_offset/$exit
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_base_plus_offset/sum_rename_req
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_word_addrgen/root_register_ack
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_base_plus_offset/sum_rename_ack
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_word_addrgen/root_register_req
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_word_addrgen/$entry
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_Update/ack
      -- CP-element group 356: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1413_Update/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(356)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(356)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(356) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr7_1405_delayed_8_0_1411_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr7_1405_delayed_8_0_1411_inst_ack_1, ack => maxPool4_CP_1841_elements(356)); -- 
    -- CP-element group 357:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	87 
    -- CP-element group 357: 	91 
    -- CP-element group 357: 	95 
    -- CP-element group 357: 	99 
    -- CP-element group 357: 	151 
    -- CP-element group 357: 	155 
    -- CP-element group 357: 	159 
    -- CP-element group 357: 	163 
    -- CP-element group 357: 	215 
    -- CP-element group 357: 	219 
    -- CP-element group 357: 	223 
    -- CP-element group 357: 	227 
    -- CP-element group 357: 	279 
    -- CP-element group 357: 	283 
    -- CP-element group 357: 	287 
    -- CP-element group 357: 	291 
    -- CP-element group 357: marked-predecessors 
    -- CP-element group 357: 	359 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_Sample/rr
      -- CP-element group 357: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_Sample/$entry
      -- CP-element group 357: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_sample_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(357)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(357)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(357) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1426_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(357), ack => CONCAT_u32_u64_1426_inst_req_0); -- 
    maxPool4_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(87) & maxPool4_CP_1841_elements(91) & maxPool4_CP_1841_elements(95) & maxPool4_CP_1841_elements(99) & maxPool4_CP_1841_elements(151) & maxPool4_CP_1841_elements(155) & maxPool4_CP_1841_elements(159) & maxPool4_CP_1841_elements(163) & maxPool4_CP_1841_elements(215) & maxPool4_CP_1841_elements(219) & maxPool4_CP_1841_elements(223) & maxPool4_CP_1841_elements(227) & maxPool4_CP_1841_elements(279) & maxPool4_CP_1841_elements(283) & maxPool4_CP_1841_elements(287) & maxPool4_CP_1841_elements(291) & maxPool4_CP_1841_elements(359);
      gj_maxPool4_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: 	363 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_Update/cr
      -- CP-element group 358: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_Update/$entry
      -- CP-element group 358: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_update_start_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(358)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(358)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(358) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1426_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(358), ack => CONCAT_u32_u64_1426_inst_req_1); -- 
    maxPool4_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(360) & maxPool4_CP_1841_elements(363);
      gj_maxPool4_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: marked-successors 
    -- CP-element group 359: 	85 
    -- CP-element group 359: 	89 
    -- CP-element group 359: 	93 
    -- CP-element group 359: 	97 
    -- CP-element group 359: 	149 
    -- CP-element group 359: 	153 
    -- CP-element group 359: 	157 
    -- CP-element group 359: 	161 
    -- CP-element group 359: 	213 
    -- CP-element group 359: 	217 
    -- CP-element group 359: 	221 
    -- CP-element group 359: 	225 
    -- CP-element group 359: 	277 
    -- CP-element group 359: 	281 
    -- CP-element group 359: 	285 
    -- CP-element group 359: 	289 
    -- CP-element group 359: 	357 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_Sample/ra
      -- CP-element group 359: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_Sample/$exit
      -- CP-element group 359: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_sample_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(359)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(359)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(359) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1426_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1426_inst_ack_0, ack => maxPool4_CP_1841_elements(359)); -- 
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	358 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_Update/ca
      -- CP-element group 360: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_Update/$exit
      -- CP-element group 360: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1426_update_completed_
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(360)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(360)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(360) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1426_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1426_inst_ack_1, ack => maxPool4_CP_1841_elements(360)); -- 
    -- CP-element group 361:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	356 
    -- CP-element group 361: 	360 
    -- CP-element group 361: 	389 
    -- CP-element group 361: marked-predecessors 
    -- CP-element group 361: 	363 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	363 
    -- CP-element group 361:  members (9) 
      -- CP-element group 361: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/$entry
      -- CP-element group 361: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_sample_start_
      -- CP-element group 361: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/ptr_deref_1415_Split/$entry
      -- CP-element group 361: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/ptr_deref_1415_Split/$exit
      -- CP-element group 361: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/ptr_deref_1415_Split/split_req
      -- CP-element group 361: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/ptr_deref_1415_Split/split_ack
      -- CP-element group 361: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/word_access_start/$entry
      -- CP-element group 361: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/word_access_start/word_0/$entry
      -- CP-element group 361: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(361)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(361)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(361) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1415_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(361), ack => ptr_deref_1415_store_0_req_0); -- 
    maxPool4_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(356) & maxPool4_CP_1841_elements(360) & maxPool4_CP_1841_elements(389) & maxPool4_CP_1841_elements(363);
      gj_maxPool4_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: marked-predecessors 
    -- CP-element group 362: 	364 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (5) 
      -- CP-element group 362: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_update_start_
      -- CP-element group 362: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Update/$entry
      -- CP-element group 362: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Update/word_access_complete/$entry
      -- CP-element group 362: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Update/word_access_complete/word_0/$entry
      -- CP-element group 362: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(362)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(362)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(362) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1415_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(362), ack => ptr_deref_1415_store_0_req_1); -- 
    maxPool4_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_1841_elements(364);
      gj_maxPool4_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	361 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	390 
    -- CP-element group 363: marked-successors 
    -- CP-element group 363: 	354 
    -- CP-element group 363: 	358 
    -- CP-element group 363: 	361 
    -- CP-element group 363:  members (5) 
      -- CP-element group 363: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_sample_completed_
      -- CP-element group 363: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/$exit
      -- CP-element group 363: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/word_access_start/$exit
      -- CP-element group 363: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/word_access_start/word_0/$exit
      -- CP-element group 363: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(363)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(363)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(363) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1415_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1415_store_0_ack_0, ack => maxPool4_CP_1841_elements(363)); -- 
    -- CP-element group 364:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	391 
    -- CP-element group 364: marked-successors 
    -- CP-element group 364: 	362 
    -- CP-element group 364:  members (5) 
      -- CP-element group 364: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_update_completed_
      -- CP-element group 364: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Update/$exit
      -- CP-element group 364: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Update/word_access_complete/$exit
      -- CP-element group 364: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Update/word_access_complete/word_0/$exit
      -- CP-element group 364: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(364)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(364)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(364) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1415_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1415_store_0_ack_1, ack => maxPool4_CP_1841_elements(364)); -- 
    -- CP-element group 365:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	369 
    -- CP-element group 365: marked-predecessors 
    -- CP-element group 365: 	370 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	370 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_sample_start_
      -- CP-element group 365: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_request/$entry
      -- CP-element group 365: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_request/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(365)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(365)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(365) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1435_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(365), ack => addr_of_1435_final_reg_req_0); -- 
    maxPool4_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(369) & maxPool4_CP_1841_elements(370);
      gj_maxPool4_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	1 
    -- CP-element group 366: marked-predecessors 
    -- CP-element group 366: 	371 
    -- CP-element group 366: 	374 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	371 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_update_start_
      -- CP-element group 366: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_complete/$entry
      -- CP-element group 366: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_complete/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(366)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(366)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(366) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1435_final_reg_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(366), ack => addr_of_1435_final_reg_req_1); -- 
    maxPool4_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(371) & maxPool4_CP_1841_elements(374);
      gj_maxPool4_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	1 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	369 
    -- CP-element group 367: 	370 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_final_index_sum_regn_update_start
      -- CP-element group 367: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_final_index_sum_regn_Update/$entry
      -- CP-element group 367: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_final_index_sum_regn_Update/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(367)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(367)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(367) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1434_index_offset_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(367), ack => array_obj_ref_1434_index_offset_req_1); -- 
    maxPool4_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(1) & maxPool4_CP_1841_elements(369) & maxPool4_CP_1841_elements(370);
      gj_maxPool4_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	1 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	391 
    -- CP-element group 368: marked-successors 
    -- CP-element group 368: 	2 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_final_index_sum_regn_sample_complete
      -- CP-element group 368: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_final_index_sum_regn_Sample/$exit
      -- CP-element group 368: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(368)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(368)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(368) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1434_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1434_index_offset_ack_0, ack => maxPool4_CP_1841_elements(368)); -- 
    -- CP-element group 369:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	365 
    -- CP-element group 369: marked-successors 
    -- CP-element group 369: 	367 
    -- CP-element group 369:  members (8) 
      -- CP-element group 369: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_root_address_calculated
      -- CP-element group 369: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_offset_calculated
      -- CP-element group 369: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_final_index_sum_regn_Update/$exit
      -- CP-element group 369: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_final_index_sum_regn_Update/ack
      -- CP-element group 369: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_base_plus_offset/$entry
      -- CP-element group 369: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_base_plus_offset/$exit
      -- CP-element group 369: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_base_plus_offset/sum_rename_req
      -- CP-element group 369: 	 assign_stmt_417_to_assign_stmt_1457/array_obj_ref_1434_base_plus_offset/sum_rename_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(369)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(369)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(369) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:array_obj_ref_1434_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1434_index_offset_ack_1, ack => maxPool4_CP_1841_elements(369)); -- 
    -- CP-element group 370:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: successors 
    -- CP-element group 370: marked-successors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: 	367 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_sample_completed_
      -- CP-element group 370: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_request/$exit
      -- CP-element group 370: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_request/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(370)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(370)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(370) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1435_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1435_final_reg_ack_0, ack => maxPool4_CP_1841_elements(370)); -- 
    -- CP-element group 371:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	366 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371: marked-successors 
    -- CP-element group 371: 	366 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_update_completed_
      -- CP-element group 371: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_complete/$exit
      -- CP-element group 371: 	 assign_stmt_417_to_assign_stmt_1457/addr_of_1435_complete/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(371)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(371)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(371) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:addr_of_1435_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1435_final_reg_ack_1, ack => maxPool4_CP_1841_elements(371)); -- 
    -- CP-element group 372:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: marked-predecessors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_sample_start_
      -- CP-element group 372: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_Sample/$entry
      -- CP-element group 372: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_Sample/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(372)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(372)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(372) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr8_1428_delayed_8_0_1437_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(372), ack => W_myptr8_1428_delayed_8_0_1437_inst_req_0); -- 
    maxPool4_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(371) & maxPool4_CP_1841_elements(374);
      gj_maxPool4_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: marked-predecessors 
    -- CP-element group 373: 	375 
    -- CP-element group 373: 	382 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_update_start_
      -- CP-element group 373: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_Update/$entry
      -- CP-element group 373: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_Update/req
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(373)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(373)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(373) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr8_1428_delayed_8_0_1437_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(373), ack => W_myptr8_1428_delayed_8_0_1437_inst_req_1); -- 
    maxPool4_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(375) & maxPool4_CP_1841_elements(382);
      gj_maxPool4_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: marked-successors 
    -- CP-element group 374: 	366 
    -- CP-element group 374: 	372 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_sample_completed_
      -- CP-element group 374: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_Sample/$exit
      -- CP-element group 374: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_Sample/ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(374)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(374)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(374) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr8_1428_delayed_8_0_1437_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr8_1428_delayed_8_0_1437_inst_ack_0, ack => maxPool4_CP_1841_elements(374)); -- 
    -- CP-element group 375:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	380 
    -- CP-element group 375: marked-successors 
    -- CP-element group 375: 	373 
    -- CP-element group 375:  members (19) 
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_update_completed_
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_Update/$exit
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/assign_stmt_1439_Update/ack
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_base_address_calculated
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_word_address_calculated
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_root_address_calculated
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_base_address_resized
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_base_addr_resize/$entry
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_base_addr_resize/$exit
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_base_addr_resize/base_resize_req
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_base_addr_resize/base_resize_ack
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_base_plus_offset/$entry
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_base_plus_offset/$exit
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_base_plus_offset/sum_rename_req
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_base_plus_offset/sum_rename_ack
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_word_addrgen/$entry
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_word_addrgen/$exit
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_word_addrgen/root_register_req
      -- CP-element group 375: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(375)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(375)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(375) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:W_myptr8_1428_delayed_8_0_1437_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr8_1428_delayed_8_0_1437_inst_ack_1, ack => maxPool4_CP_1841_elements(375)); -- 
    -- CP-element group 376:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	103 
    -- CP-element group 376: 	107 
    -- CP-element group 376: 	111 
    -- CP-element group 376: 	115 
    -- CP-element group 376: 	167 
    -- CP-element group 376: 	171 
    -- CP-element group 376: 	175 
    -- CP-element group 376: 	179 
    -- CP-element group 376: 	231 
    -- CP-element group 376: 	235 
    -- CP-element group 376: 	239 
    -- CP-element group 376: 	243 
    -- CP-element group 376: 	295 
    -- CP-element group 376: 	299 
    -- CP-element group 376: 	303 
    -- CP-element group 376: 	307 
    -- CP-element group 376: marked-predecessors 
    -- CP-element group 376: 	378 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	378 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_sample_start_
      -- CP-element group 376: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_Sample/$entry
      -- CP-element group 376: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(376)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(376)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(376) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1452_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(376), ack => CONCAT_u32_u64_1452_inst_req_0); -- 
    maxPool4_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(103) & maxPool4_CP_1841_elements(107) & maxPool4_CP_1841_elements(111) & maxPool4_CP_1841_elements(115) & maxPool4_CP_1841_elements(167) & maxPool4_CP_1841_elements(171) & maxPool4_CP_1841_elements(175) & maxPool4_CP_1841_elements(179) & maxPool4_CP_1841_elements(231) & maxPool4_CP_1841_elements(235) & maxPool4_CP_1841_elements(239) & maxPool4_CP_1841_elements(243) & maxPool4_CP_1841_elements(295) & maxPool4_CP_1841_elements(299) & maxPool4_CP_1841_elements(303) & maxPool4_CP_1841_elements(307) & maxPool4_CP_1841_elements(378);
      gj_maxPool4_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: marked-predecessors 
    -- CP-element group 377: 	379 
    -- CP-element group 377: 	382 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_update_start_
      -- CP-element group 377: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_Update/$entry
      -- CP-element group 377: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(377)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(377)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(377) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1452_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(377), ack => CONCAT_u32_u64_1452_inst_req_1); -- 
    maxPool4_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(379) & maxPool4_CP_1841_elements(382);
      gj_maxPool4_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	376 
    -- CP-element group 378: successors 
    -- CP-element group 378: marked-successors 
    -- CP-element group 378: 	101 
    -- CP-element group 378: 	105 
    -- CP-element group 378: 	109 
    -- CP-element group 378: 	113 
    -- CP-element group 378: 	165 
    -- CP-element group 378: 	169 
    -- CP-element group 378: 	173 
    -- CP-element group 378: 	177 
    -- CP-element group 378: 	229 
    -- CP-element group 378: 	233 
    -- CP-element group 378: 	237 
    -- CP-element group 378: 	241 
    -- CP-element group 378: 	293 
    -- CP-element group 378: 	297 
    -- CP-element group 378: 	301 
    -- CP-element group 378: 	305 
    -- CP-element group 378: 	376 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_sample_completed_
      -- CP-element group 378: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_Sample/$exit
      -- CP-element group 378: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(378)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(378)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(378) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1452_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1452_inst_ack_0, ack => maxPool4_CP_1841_elements(378)); -- 
    -- CP-element group 379:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379: marked-successors 
    -- CP-element group 379: 	377 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_update_completed_
      -- CP-element group 379: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_Update/$exit
      -- CP-element group 379: 	 assign_stmt_417_to_assign_stmt_1457/CONCAT_u32_u64_1452_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(379)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(379)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(379) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:CONCAT_u32_u64_1452_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1452_inst_ack_1, ack => maxPool4_CP_1841_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	375 
    -- CP-element group 380: 	379 
    -- CP-element group 380: 	390 
    -- CP-element group 380: marked-predecessors 
    -- CP-element group 380: 	382 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (9) 
      -- CP-element group 380: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_sample_start_
      -- CP-element group 380: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/$entry
      -- CP-element group 380: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/ptr_deref_1441_Split/$entry
      -- CP-element group 380: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/ptr_deref_1441_Split/$exit
      -- CP-element group 380: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/ptr_deref_1441_Split/split_req
      -- CP-element group 380: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/ptr_deref_1441_Split/split_ack
      -- CP-element group 380: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/word_access_start/$entry
      -- CP-element group 380: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/word_access_start/word_0/$entry
      -- CP-element group 380: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(380)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(380)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(380) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1441_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(380), ack => ptr_deref_1441_store_0_req_0); -- 
    maxPool4_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(375) & maxPool4_CP_1841_elements(379) & maxPool4_CP_1841_elements(390) & maxPool4_CP_1841_elements(382);
      gj_maxPool4_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: marked-predecessors 
    -- CP-element group 381: 	383 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	383 
    -- CP-element group 381:  members (5) 
      -- CP-element group 381: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_update_start_
      -- CP-element group 381: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Update/$entry
      -- CP-element group 381: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Update/word_access_complete/$entry
      -- CP-element group 381: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Update/word_access_complete/word_0/$entry
      -- CP-element group 381: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(381)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(381)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(381) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1441_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(381), ack => ptr_deref_1441_store_0_req_1); -- 
    maxPool4_cp_element_group_381: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_381"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_1841_elements(383);
      gj_maxPool4_cp_element_group_381 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(381), clk => clk, reset => reset); --
    end block;
    -- CP-element group 382:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	391 
    -- CP-element group 382: marked-successors 
    -- CP-element group 382: 	323 
    -- CP-element group 382: 	373 
    -- CP-element group 382: 	377 
    -- CP-element group 382: 	380 
    -- CP-element group 382:  members (6) 
      -- CP-element group 382: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_sample_completed_
      -- CP-element group 382: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/$exit
      -- CP-element group 382: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/word_access_start/$exit
      -- CP-element group 382: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/word_access_start/word_0/$exit
      -- CP-element group 382: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Sample/word_access_start/word_0/ra
      -- CP-element group 382: 	 assign_stmt_417_to_assign_stmt_1457/ring_reenable_memory_space_0
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(382)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(382)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(382) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1441_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1441_store_0_ack_0, ack => maxPool4_CP_1841_elements(382)); -- 
    -- CP-element group 383:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	381 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	391 
    -- CP-element group 383: marked-successors 
    -- CP-element group 383: 	381 
    -- CP-element group 383:  members (5) 
      -- CP-element group 383: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_update_completed_
      -- CP-element group 383: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Update/$exit
      -- CP-element group 383: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Update/word_access_complete/$exit
      -- CP-element group 383: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Update/word_access_complete/word_0/$exit
      -- CP-element group 383: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1441_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(383)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(383)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(383) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:ptr_deref_1441_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1441_store_0_ack_1, ack => maxPool4_CP_1841_elements(383)); -- 
    -- CP-element group 384:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	55 
    -- CP-element group 384: 	119 
    -- CP-element group 384: 	183 
    -- CP-element group 384: 	247 
    -- CP-element group 384: marked-predecessors 
    -- CP-element group 384: 	386 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	386 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_sample_start_
      -- CP-element group 384: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_Sample/$entry
      -- CP-element group 384: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_Sample/rr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(384)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(384)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(384) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:type_cast_1456_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(384), ack => type_cast_1456_inst_req_0); -- 
    maxPool4_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(55) & maxPool4_CP_1841_elements(119) & maxPool4_CP_1841_elements(183) & maxPool4_CP_1841_elements(247) & maxPool4_CP_1841_elements(386);
      gj_maxPool4_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	7 
    -- CP-element group 385: marked-predecessors 
    -- CP-element group 385: 	387 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	387 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_update_start_
      -- CP-element group 385: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_Update/$entry
      -- CP-element group 385: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_Update/cr
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(385)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(385)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(385) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:type_cast_1456_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_1841_elements(385), ack => type_cast_1456_inst_req_1); -- 
    maxPool4_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(7) & maxPool4_CP_1841_elements(387);
      gj_maxPool4_cp_element_group_385 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	384 
    -- CP-element group 386: successors 
    -- CP-element group 386: marked-successors 
    -- CP-element group 386: 	53 
    -- CP-element group 386: 	117 
    -- CP-element group 386: 	181 
    -- CP-element group 386: 	245 
    -- CP-element group 386: 	384 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_sample_completed_
      -- CP-element group 386: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_Sample/$exit
      -- CP-element group 386: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_Sample/ra
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(386)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(386)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(386) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:type_cast_1456_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1456_inst_ack_0, ack => maxPool4_CP_1841_elements(386)); -- 
    -- CP-element group 387:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	385 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	391 
    -- CP-element group 387: marked-successors 
    -- CP-element group 387: 	385 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_update_completed_
      -- CP-element group 387: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_Update/$exit
      -- CP-element group 387: 	 assign_stmt_417_to_assign_stmt_1457/type_cast_1456_Update/ca
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(387)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(387)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(387) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:type_cast_1456_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1456_inst_ack_1, ack => maxPool4_CP_1841_elements(387)); -- 
    -- CP-element group 388:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	325 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	342 
    -- CP-element group 388:  members (1) 
      -- CP-element group 388: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1363_ptr_deref_1389_delay
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(388)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(388)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(388) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool4_CP_1841_elements(388) is a control-delay.
    cp_element_388_delay: control_delay_element  generic map(name => " 388_delay", delay_value => 1)  port map(req => maxPool4_CP_1841_elements(325), ack => maxPool4_CP_1841_elements(388), clk => clk, reset =>reset);
    -- CP-element group 389:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	344 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	361 
    -- CP-element group 389:  members (1) 
      -- CP-element group 389: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1389_ptr_deref_1415_delay
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(389)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(389)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(389) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool4_CP_1841_elements(389) is a control-delay.
    cp_element_389_delay: control_delay_element  generic map(name => " 389_delay", delay_value => 1)  port map(req => maxPool4_CP_1841_elements(344), ack => maxPool4_CP_1841_elements(389), clk => clk, reset =>reset);
    -- CP-element group 390:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	363 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	380 
    -- CP-element group 390:  members (1) 
      -- CP-element group 390: 	 assign_stmt_417_to_assign_stmt_1457/ptr_deref_1415_ptr_deref_1441_delay
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(390)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(390)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(390) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group maxPool4_CP_1841_elements(390) is a control-delay.
    cp_element_390_delay: control_delay_element  generic map(name => " 390_delay", delay_value => 1)  port map(req => maxPool4_CP_1841_elements(363), ack => maxPool4_CP_1841_elements(390), clk => clk, reset =>reset);
    -- CP-element group 391:  join  transition  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	11 
    -- CP-element group 391: 	18 
    -- CP-element group 391: 	25 
    -- CP-element group 391: 	32 
    -- CP-element group 391: 	311 
    -- CP-element group 391: 	326 
    -- CP-element group 391: 	330 
    -- CP-element group 391: 	345 
    -- CP-element group 391: 	349 
    -- CP-element group 391: 	364 
    -- CP-element group 391: 	368 
    -- CP-element group 391: 	382 
    -- CP-element group 391: 	383 
    -- CP-element group 391: 	387 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	398 
    -- CP-element group 391:  members (1) 
      -- CP-element group 391: 	 assign_stmt_417_to_assign_stmt_1457/$exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(391)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(391)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(391) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= maxPool4_CP_1841_elements(11) & maxPool4_CP_1841_elements(18) & maxPool4_CP_1841_elements(25) & maxPool4_CP_1841_elements(32) & maxPool4_CP_1841_elements(311) & maxPool4_CP_1841_elements(326) & maxPool4_CP_1841_elements(330) & maxPool4_CP_1841_elements(345) & maxPool4_CP_1841_elements(349) & maxPool4_CP_1841_elements(364) & maxPool4_CP_1841_elements(368) & maxPool4_CP_1841_elements(382) & maxPool4_CP_1841_elements(383) & maxPool4_CP_1841_elements(387);
      gj_maxPool4_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_1841_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  place  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	2 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (1) 
      -- CP-element group 392: 	 addr_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(392)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(392)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(392) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_CP_1841_elements(392) <= maxPool4_CP_1841_elements(2);
    -- CP-element group 393:  place  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	3 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (1) 
      -- CP-element group 393: 	 addr1_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(393)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(393)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(393) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_CP_1841_elements(393) <= maxPool4_CP_1841_elements(3);
    -- CP-element group 394:  place  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	4 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (1) 
      -- CP-element group 394: 	 addr2_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(394)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(394)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(394) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_CP_1841_elements(394) <= maxPool4_CP_1841_elements(4);
    -- CP-element group 395:  place  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	5 
    -- CP-element group 395: successors 
    -- CP-element group 395:  members (1) 
      -- CP-element group 395: 	 addr3_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(395)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(395)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(395) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_CP_1841_elements(395) <= maxPool4_CP_1841_elements(5);
    -- CP-element group 396:  place  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	6 
    -- CP-element group 396: successors 
    -- CP-element group 396:  members (1) 
      -- CP-element group 396: 	 addr4_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(396)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(396)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(396) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_CP_1841_elements(396) <= maxPool4_CP_1841_elements(6);
    -- CP-element group 397:  place  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	7 
    -- CP-element group 397:  members (1) 
      -- CP-element group 397: 	 output_update_enable
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(397)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(397)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(397) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 398:  transition  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	391 
    -- CP-element group 398: successors 
    -- CP-element group 398:  members (1) 
      -- CP-element group 398: 	 $exit
      -- 
    -- logger for CP element group maxPool4_CP_1841_elements(398)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and maxPool4_CP_1841_elements(398)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:maxPool4:CP:maxPool4_CP_1841_elements(398) fired."); 
        -- 
      end if; --
    end process; 
    maxPool4_CP_1841_elements(398) <= maxPool4_CP_1841_elements(391);
    --  hookup: inputs to control-path 
    maxPool4_CP_1841_elements(397) <= output_update_enable;
    -- hookup: output from control-path 
    addr_update_enable <= maxPool4_CP_1841_elements(392);
    addr1_update_enable <= maxPool4_CP_1841_elements(393);
    addr2_update_enable <= maxPool4_CP_1841_elements(394);
    addr3_update_enable <= maxPool4_CP_1841_elements(395);
    addr4_update_enable <= maxPool4_CP_1841_elements(396);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1381_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1381_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1381_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1407_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1407_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1407_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1433_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1433_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1433_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1368_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1373_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1394_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1399_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1420_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1425_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1446_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1451_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_1374_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1400_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1426_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1452_wire : std_logic_vector(63 downto 0);
    signal R_addr1_414_resized : std_logic_vector(13 downto 0);
    signal R_addr1_414_scaled : std_logic_vector(13 downto 0);
    signal R_addr2_421_resized : std_logic_vector(13 downto 0);
    signal R_addr2_421_scaled : std_logic_vector(13 downto 0);
    signal R_addr3_428_resized : std_logic_vector(13 downto 0);
    signal R_addr3_428_scaled : std_logic_vector(13 downto 0);
    signal R_addr4_435_resized : std_logic_vector(13 downto 0);
    signal R_addr4_435_scaled : std_logic_vector(13 downto 0);
    signal R_addr_1355_resized : std_logic_vector(13 downto 0);
    signal R_addr_1355_scaled : std_logic_vector(13 downto 0);
    signal SGT_i16_u1_1003_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1011_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1019_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1027_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1035_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1043_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1051_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1059_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1067_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1075_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1083_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1091_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1099_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1107_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1115_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1123_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1131_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1139_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1147_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1155_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1163_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1171_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1179_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1187_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1195_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1203_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1211_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1219_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1227_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1235_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1243_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1251_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1259_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1267_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1275_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1283_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1291_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1299_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1307_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1315_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1323_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1331_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1339_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1347_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_971_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_979_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_987_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_995_wire : std_logic_vector(0 downto 0);
    signal a110_751 : std_logic_vector(15 downto 0);
    signal a111_755 : std_logic_vector(15 downto 0);
    signal a112_759 : std_logic_vector(15 downto 0);
    signal a113_763 : std_logic_vector(15 downto 0);
    signal a114_767 : std_logic_vector(15 downto 0);
    signal a115_771 : std_logic_vector(15 downto 0);
    signal a116_775 : std_logic_vector(15 downto 0);
    signal a11_715 : std_logic_vector(15 downto 0);
    signal a12_719 : std_logic_vector(15 downto 0);
    signal a13_723 : std_logic_vector(15 downto 0);
    signal a14_727 : std_logic_vector(15 downto 0);
    signal a15_731 : std_logic_vector(15 downto 0);
    signal a16_735 : std_logic_vector(15 downto 0);
    signal a17_739 : std_logic_vector(15 downto 0);
    signal a18_743 : std_logic_vector(15 downto 0);
    signal a19_747 : std_logic_vector(15 downto 0);
    signal a210_815 : std_logic_vector(15 downto 0);
    signal a211_819 : std_logic_vector(15 downto 0);
    signal a212_823 : std_logic_vector(15 downto 0);
    signal a213_827 : std_logic_vector(15 downto 0);
    signal a214_831 : std_logic_vector(15 downto 0);
    signal a215_835 : std_logic_vector(15 downto 0);
    signal a216_839 : std_logic_vector(15 downto 0);
    signal a21_779 : std_logic_vector(15 downto 0);
    signal a22_783 : std_logic_vector(15 downto 0);
    signal a23_787 : std_logic_vector(15 downto 0);
    signal a24_791 : std_logic_vector(15 downto 0);
    signal a25_795 : std_logic_vector(15 downto 0);
    signal a26_799 : std_logic_vector(15 downto 0);
    signal a27_803 : std_logic_vector(15 downto 0);
    signal a28_807 : std_logic_vector(15 downto 0);
    signal a29_811 : std_logic_vector(15 downto 0);
    signal a310_879 : std_logic_vector(15 downto 0);
    signal a311_883 : std_logic_vector(15 downto 0);
    signal a312_887 : std_logic_vector(15 downto 0);
    signal a313_891 : std_logic_vector(15 downto 0);
    signal a314_895 : std_logic_vector(15 downto 0);
    signal a315_899 : std_logic_vector(15 downto 0);
    signal a316_903 : std_logic_vector(15 downto 0);
    signal a31_843 : std_logic_vector(15 downto 0);
    signal a32_847 : std_logic_vector(15 downto 0);
    signal a33_851 : std_logic_vector(15 downto 0);
    signal a34_855 : std_logic_vector(15 downto 0);
    signal a35_859 : std_logic_vector(15 downto 0);
    signal a36_863 : std_logic_vector(15 downto 0);
    signal a37_867 : std_logic_vector(15 downto 0);
    signal a38_871 : std_logic_vector(15 downto 0);
    signal a39_875 : std_logic_vector(15 downto 0);
    signal a410_943 : std_logic_vector(15 downto 0);
    signal a411_947 : std_logic_vector(15 downto 0);
    signal a412_951 : std_logic_vector(15 downto 0);
    signal a413_955 : std_logic_vector(15 downto 0);
    signal a414_959 : std_logic_vector(15 downto 0);
    signal a415_963 : std_logic_vector(15 downto 0);
    signal a416_967 : std_logic_vector(15 downto 0);
    signal a41_907 : std_logic_vector(15 downto 0);
    signal a42_911 : std_logic_vector(15 downto 0);
    signal a43_915 : std_logic_vector(15 downto 0);
    signal a44_919 : std_logic_vector(15 downto 0);
    signal a45_923 : std_logic_vector(15 downto 0);
    signal a46_927 : std_logic_vector(15 downto 0);
    signal a47_931 : std_logic_vector(15 downto 0);
    signal a48_935 : std_logic_vector(15 downto 0);
    signal a49_939 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1356_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1356_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1356_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1356_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1356_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1356_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1382_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1382_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1382_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1382_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1382_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1382_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1434_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1434_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1434_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1434_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1434_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1434_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_422_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_422_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_422_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_422_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_422_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_422_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_429_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_429_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_429_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_429_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_429_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_429_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_436_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_436_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_436_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_436_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_436_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_436_root_address : std_logic_vector(13 downto 0);
    signal c1_442 : std_logic_vector(255 downto 0);
    signal c2_446 : std_logic_vector(255 downto 0);
    signal c3_450 : std_logic_vector(255 downto 0);
    signal c4_454 : std_logic_vector(255 downto 0);
    signal konst_1380_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1406_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1432_wire_constant : std_logic_vector(31 downto 0);
    signal myptr1_417 : std_logic_vector(31 downto 0);
    signal myptr2_424 : std_logic_vector(31 downto 0);
    signal myptr3_431 : std_logic_vector(31 downto 0);
    signal myptr4_438 : std_logic_vector(31 downto 0);
    signal myptr5_1358 : std_logic_vector(31 downto 0);
    signal myptr5_1359_delayed_8_0_1361 : std_logic_vector(31 downto 0);
    signal myptr6_1382_delayed_8_0_1387 : std_logic_vector(31 downto 0);
    signal myptr6_1384 : std_logic_vector(31 downto 0);
    signal myptr7_1405_delayed_8_0_1413 : std_logic_vector(31 downto 0);
    signal myptr7_1410 : std_logic_vector(31 downto 0);
    signal myptr8_1428_delayed_8_0_1439 : std_logic_vector(31 downto 0);
    signal myptr8_1436 : std_logic_vector(31 downto 0);
    signal out10_1207 : std_logic_vector(15 downto 0);
    signal out11_1231 : std_logic_vector(15 downto 0);
    signal out12_1255 : std_logic_vector(15 downto 0);
    signal out13_1279 : std_logic_vector(15 downto 0);
    signal out14_1303 : std_logic_vector(15 downto 0);
    signal out15_1327 : std_logic_vector(15 downto 0);
    signal out16_1351 : std_logic_vector(15 downto 0);
    signal out1_991 : std_logic_vector(15 downto 0);
    signal out2_1015 : std_logic_vector(15 downto 0);
    signal out3_1039 : std_logic_vector(15 downto 0);
    signal out4_1063 : std_logic_vector(15 downto 0);
    signal out5_1087 : std_logic_vector(15 downto 0);
    signal out6_1111 : std_logic_vector(15 downto 0);
    signal out7_1135 : std_logic_vector(15 downto 0);
    signal out8_1159 : std_logic_vector(15 downto 0);
    signal out9_1183 : std_logic_vector(15 downto 0);
    signal ptr_deref_1363_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1363_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1363_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1363_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1363_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1363_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1389_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1389_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1389_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1389_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1389_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1389_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1415_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1415_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1415_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1415_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1415_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1415_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1441_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1441_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1441_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1441_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1441_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1441_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_441_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_441_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_441_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_441_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_441_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_445_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_445_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_445_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_445_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_445_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_449_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_449_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_449_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_449_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_449_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_453_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_453_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_453_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_453_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_453_word_offset_0 : std_logic_vector(13 downto 0);
    signal sliced_v110_494 : std_logic_vector(15 downto 0);
    signal sliced_v111_498 : std_logic_vector(15 downto 0);
    signal sliced_v112_502 : std_logic_vector(15 downto 0);
    signal sliced_v113_506 : std_logic_vector(15 downto 0);
    signal sliced_v114_510 : std_logic_vector(15 downto 0);
    signal sliced_v115_514 : std_logic_vector(15 downto 0);
    signal sliced_v116_518 : std_logic_vector(15 downto 0);
    signal sliced_v11_458 : std_logic_vector(15 downto 0);
    signal sliced_v12_462 : std_logic_vector(15 downto 0);
    signal sliced_v13_466 : std_logic_vector(15 downto 0);
    signal sliced_v14_470 : std_logic_vector(15 downto 0);
    signal sliced_v15_474 : std_logic_vector(15 downto 0);
    signal sliced_v16_478 : std_logic_vector(15 downto 0);
    signal sliced_v17_482 : std_logic_vector(15 downto 0);
    signal sliced_v18_486 : std_logic_vector(15 downto 0);
    signal sliced_v19_490 : std_logic_vector(15 downto 0);
    signal sliced_v210_558 : std_logic_vector(15 downto 0);
    signal sliced_v211_562 : std_logic_vector(15 downto 0);
    signal sliced_v212_566 : std_logic_vector(15 downto 0);
    signal sliced_v213_570 : std_logic_vector(15 downto 0);
    signal sliced_v214_574 : std_logic_vector(15 downto 0);
    signal sliced_v215_578 : std_logic_vector(15 downto 0);
    signal sliced_v216_582 : std_logic_vector(15 downto 0);
    signal sliced_v21_522 : std_logic_vector(15 downto 0);
    signal sliced_v22_526 : std_logic_vector(15 downto 0);
    signal sliced_v23_530 : std_logic_vector(15 downto 0);
    signal sliced_v24_534 : std_logic_vector(15 downto 0);
    signal sliced_v25_538 : std_logic_vector(15 downto 0);
    signal sliced_v26_542 : std_logic_vector(15 downto 0);
    signal sliced_v27_546 : std_logic_vector(15 downto 0);
    signal sliced_v28_550 : std_logic_vector(15 downto 0);
    signal sliced_v29_554 : std_logic_vector(15 downto 0);
    signal sliced_v310_622 : std_logic_vector(15 downto 0);
    signal sliced_v311_626 : std_logic_vector(15 downto 0);
    signal sliced_v312_630 : std_logic_vector(15 downto 0);
    signal sliced_v313_634 : std_logic_vector(15 downto 0);
    signal sliced_v314_638 : std_logic_vector(15 downto 0);
    signal sliced_v315_642 : std_logic_vector(15 downto 0);
    signal sliced_v316_646 : std_logic_vector(15 downto 0);
    signal sliced_v31_586 : std_logic_vector(15 downto 0);
    signal sliced_v32_590 : std_logic_vector(15 downto 0);
    signal sliced_v33_594 : std_logic_vector(15 downto 0);
    signal sliced_v34_598 : std_logic_vector(15 downto 0);
    signal sliced_v35_602 : std_logic_vector(15 downto 0);
    signal sliced_v36_606 : std_logic_vector(15 downto 0);
    signal sliced_v37_610 : std_logic_vector(15 downto 0);
    signal sliced_v38_614 : std_logic_vector(15 downto 0);
    signal sliced_v39_618 : std_logic_vector(15 downto 0);
    signal sliced_v410_686 : std_logic_vector(15 downto 0);
    signal sliced_v411_690 : std_logic_vector(15 downto 0);
    signal sliced_v412_694 : std_logic_vector(15 downto 0);
    signal sliced_v413_698 : std_logic_vector(15 downto 0);
    signal sliced_v414_702 : std_logic_vector(15 downto 0);
    signal sliced_v415_706 : std_logic_vector(15 downto 0);
    signal sliced_v416_710 : std_logic_vector(15 downto 0);
    signal sliced_v41_650 : std_logic_vector(15 downto 0);
    signal sliced_v42_654 : std_logic_vector(15 downto 0);
    signal sliced_v43_658 : std_logic_vector(15 downto 0);
    signal sliced_v44_662 : std_logic_vector(15 downto 0);
    signal sliced_v45_666 : std_logic_vector(15 downto 0);
    signal sliced_v46_670 : std_logic_vector(15 downto 0);
    signal sliced_v47_674 : std_logic_vector(15 downto 0);
    signal sliced_v48_678 : std_logic_vector(15 downto 0);
    signal sliced_v49_682 : std_logic_vector(15 downto 0);
    signal t101_1191 : std_logic_vector(15 downto 0);
    signal t102_1199 : std_logic_vector(15 downto 0);
    signal t111_1215 : std_logic_vector(15 downto 0);
    signal t112_1223 : std_logic_vector(15 downto 0);
    signal t11_975 : std_logic_vector(15 downto 0);
    signal t121_1239 : std_logic_vector(15 downto 0);
    signal t122_1247 : std_logic_vector(15 downto 0);
    signal t12_983 : std_logic_vector(15 downto 0);
    signal t131_1263 : std_logic_vector(15 downto 0);
    signal t132_1271 : std_logic_vector(15 downto 0);
    signal t141_1287 : std_logic_vector(15 downto 0);
    signal t142_1295 : std_logic_vector(15 downto 0);
    signal t151_1311 : std_logic_vector(15 downto 0);
    signal t152_1319 : std_logic_vector(15 downto 0);
    signal t161_1335 : std_logic_vector(15 downto 0);
    signal t162_1343 : std_logic_vector(15 downto 0);
    signal t21_999 : std_logic_vector(15 downto 0);
    signal t22_1007 : std_logic_vector(15 downto 0);
    signal t31_1023 : std_logic_vector(15 downto 0);
    signal t32_1031 : std_logic_vector(15 downto 0);
    signal t41_1047 : std_logic_vector(15 downto 0);
    signal t42_1055 : std_logic_vector(15 downto 0);
    signal t51_1071 : std_logic_vector(15 downto 0);
    signal t52_1079 : std_logic_vector(15 downto 0);
    signal t61_1095 : std_logic_vector(15 downto 0);
    signal t62_1103 : std_logic_vector(15 downto 0);
    signal t71_1119 : std_logic_vector(15 downto 0);
    signal t72_1127 : std_logic_vector(15 downto 0);
    signal t81_1143 : std_logic_vector(15 downto 0);
    signal t82_1151 : std_logic_vector(15 downto 0);
    signal t91_1167 : std_logic_vector(15 downto 0);
    signal t92_1175 : std_logic_vector(15 downto 0);
    signal type_cast_1365_wire : std_logic_vector(15 downto 0);
    signal type_cast_1367_wire : std_logic_vector(15 downto 0);
    signal type_cast_1370_wire : std_logic_vector(15 downto 0);
    signal type_cast_1372_wire : std_logic_vector(15 downto 0);
    signal type_cast_1391_wire : std_logic_vector(15 downto 0);
    signal type_cast_1393_wire : std_logic_vector(15 downto 0);
    signal type_cast_1396_wire : std_logic_vector(15 downto 0);
    signal type_cast_1398_wire : std_logic_vector(15 downto 0);
    signal type_cast_1417_wire : std_logic_vector(15 downto 0);
    signal type_cast_1419_wire : std_logic_vector(15 downto 0);
    signal type_cast_1422_wire : std_logic_vector(15 downto 0);
    signal type_cast_1424_wire : std_logic_vector(15 downto 0);
    signal type_cast_1443_wire : std_logic_vector(15 downto 0);
    signal type_cast_1445_wire : std_logic_vector(15 downto 0);
    signal type_cast_1448_wire : std_logic_vector(15 downto 0);
    signal type_cast_1450_wire : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1356_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1356_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1356_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1356_resized_base_address <= "00000000000000";
    array_obj_ref_1382_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1382_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1382_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1382_resized_base_address <= "00000000000000";
    array_obj_ref_1408_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1408_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1408_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1408_resized_base_address <= "00000000000000";
    array_obj_ref_1434_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1434_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1434_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1434_resized_base_address <= "00000000000000";
    array_obj_ref_415_constant_part_of_offset <= "00000000000000";
    array_obj_ref_415_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_415_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_415_resized_base_address <= "00000000000000";
    array_obj_ref_422_constant_part_of_offset <= "00000000000000";
    array_obj_ref_422_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_422_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_422_resized_base_address <= "00000000000000";
    array_obj_ref_429_constant_part_of_offset <= "00000000000000";
    array_obj_ref_429_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_429_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_429_resized_base_address <= "00000000000000";
    array_obj_ref_436_constant_part_of_offset <= "00000000000000";
    array_obj_ref_436_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_436_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_436_resized_base_address <= "00000000000000";
    konst_1380_wire_constant <= "00000000000000000000000000000001";
    konst_1406_wire_constant <= "00000000000000000000000000000010";
    konst_1432_wire_constant <= "00000000000000000000000000000011";
    ptr_deref_1363_word_offset_0 <= "00000000000000";
    ptr_deref_1389_word_offset_0 <= "00000000000000";
    ptr_deref_1415_word_offset_0 <= "00000000000000";
    ptr_deref_1441_word_offset_0 <= "00000000000000";
    ptr_deref_441_word_offset_0 <= "00000000000000";
    ptr_deref_445_word_offset_0 <= "00000000000000";
    ptr_deref_449_word_offset_0 <= "00000000000000";
    ptr_deref_453_word_offset_0 <= "00000000000000";
    -- logger for split-operator MUX_1006_inst flow-through 
    process(t22_1007) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1006_inst:flowthrough inputs: " & " SGT_i16_u1_1003_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1003_wire) & " a32_847 = "& Convert_SLV_To_Hex_String(a32_847) & " a42_911 = "& Convert_SLV_To_Hex_String(a42_911) & " outputs:" & " t22_1007= "  & Convert_SLV_To_Hex_String(t22_1007));
      --
    end process; 
    -- flow-through select operator MUX_1006_inst
    t22_1007 <= a32_847 when (SGT_i16_u1_1003_wire(0) /=  '0') else a42_911;
    -- logger for split-operator MUX_1014_inst flow-through 
    process(out2_1015) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1014_inst:flowthrough inputs: " & " SGT_i16_u1_1011_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1011_wire) & " t21_999 = "& Convert_SLV_To_Hex_String(t21_999) & " t22_1007 = "& Convert_SLV_To_Hex_String(t22_1007) & " outputs:" & " out2_1015= "  & Convert_SLV_To_Hex_String(out2_1015));
      --
    end process; 
    -- flow-through select operator MUX_1014_inst
    out2_1015 <= t21_999 when (SGT_i16_u1_1011_wire(0) /=  '0') else t22_1007;
    -- logger for split-operator MUX_1022_inst flow-through 
    process(t31_1023) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1022_inst:flowthrough inputs: " & " SGT_i16_u1_1019_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1019_wire) & " a13_723 = "& Convert_SLV_To_Hex_String(a13_723) & " a23_787 = "& Convert_SLV_To_Hex_String(a23_787) & " outputs:" & " t31_1023= "  & Convert_SLV_To_Hex_String(t31_1023));
      --
    end process; 
    -- flow-through select operator MUX_1022_inst
    t31_1023 <= a13_723 when (SGT_i16_u1_1019_wire(0) /=  '0') else a23_787;
    -- logger for split-operator MUX_1030_inst flow-through 
    process(t32_1031) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1030_inst:flowthrough inputs: " & " SGT_i16_u1_1027_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1027_wire) & " a33_851 = "& Convert_SLV_To_Hex_String(a33_851) & " a43_915 = "& Convert_SLV_To_Hex_String(a43_915) & " outputs:" & " t32_1031= "  & Convert_SLV_To_Hex_String(t32_1031));
      --
    end process; 
    -- flow-through select operator MUX_1030_inst
    t32_1031 <= a33_851 when (SGT_i16_u1_1027_wire(0) /=  '0') else a43_915;
    -- logger for split-operator MUX_1038_inst flow-through 
    process(out3_1039) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1038_inst:flowthrough inputs: " & " SGT_i16_u1_1035_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1035_wire) & " t31_1023 = "& Convert_SLV_To_Hex_String(t31_1023) & " t32_1031 = "& Convert_SLV_To_Hex_String(t32_1031) & " outputs:" & " out3_1039= "  & Convert_SLV_To_Hex_String(out3_1039));
      --
    end process; 
    -- flow-through select operator MUX_1038_inst
    out3_1039 <= t31_1023 when (SGT_i16_u1_1035_wire(0) /=  '0') else t32_1031;
    -- logger for split-operator MUX_1046_inst flow-through 
    process(t41_1047) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1046_inst:flowthrough inputs: " & " SGT_i16_u1_1043_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1043_wire) & " a14_727 = "& Convert_SLV_To_Hex_String(a14_727) & " a24_791 = "& Convert_SLV_To_Hex_String(a24_791) & " outputs:" & " t41_1047= "  & Convert_SLV_To_Hex_String(t41_1047));
      --
    end process; 
    -- flow-through select operator MUX_1046_inst
    t41_1047 <= a14_727 when (SGT_i16_u1_1043_wire(0) /=  '0') else a24_791;
    -- logger for split-operator MUX_1054_inst flow-through 
    process(t42_1055) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1054_inst:flowthrough inputs: " & " SGT_i16_u1_1051_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1051_wire) & " a34_855 = "& Convert_SLV_To_Hex_String(a34_855) & " a44_919 = "& Convert_SLV_To_Hex_String(a44_919) & " outputs:" & " t42_1055= "  & Convert_SLV_To_Hex_String(t42_1055));
      --
    end process; 
    -- flow-through select operator MUX_1054_inst
    t42_1055 <= a34_855 when (SGT_i16_u1_1051_wire(0) /=  '0') else a44_919;
    -- logger for split-operator MUX_1062_inst flow-through 
    process(out4_1063) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1062_inst:flowthrough inputs: " & " SGT_i16_u1_1059_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1059_wire) & " t41_1047 = "& Convert_SLV_To_Hex_String(t41_1047) & " t42_1055 = "& Convert_SLV_To_Hex_String(t42_1055) & " outputs:" & " out4_1063= "  & Convert_SLV_To_Hex_String(out4_1063));
      --
    end process; 
    -- flow-through select operator MUX_1062_inst
    out4_1063 <= t41_1047 when (SGT_i16_u1_1059_wire(0) /=  '0') else t42_1055;
    -- logger for split-operator MUX_1070_inst flow-through 
    process(t51_1071) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1070_inst:flowthrough inputs: " & " SGT_i16_u1_1067_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1067_wire) & " a15_731 = "& Convert_SLV_To_Hex_String(a15_731) & " a25_795 = "& Convert_SLV_To_Hex_String(a25_795) & " outputs:" & " t51_1071= "  & Convert_SLV_To_Hex_String(t51_1071));
      --
    end process; 
    -- flow-through select operator MUX_1070_inst
    t51_1071 <= a15_731 when (SGT_i16_u1_1067_wire(0) /=  '0') else a25_795;
    -- logger for split-operator MUX_1078_inst flow-through 
    process(t52_1079) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1078_inst:flowthrough inputs: " & " SGT_i16_u1_1075_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1075_wire) & " a35_859 = "& Convert_SLV_To_Hex_String(a35_859) & " a45_923 = "& Convert_SLV_To_Hex_String(a45_923) & " outputs:" & " t52_1079= "  & Convert_SLV_To_Hex_String(t52_1079));
      --
    end process; 
    -- flow-through select operator MUX_1078_inst
    t52_1079 <= a35_859 when (SGT_i16_u1_1075_wire(0) /=  '0') else a45_923;
    -- logger for split-operator MUX_1086_inst flow-through 
    process(out5_1087) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1086_inst:flowthrough inputs: " & " SGT_i16_u1_1083_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1083_wire) & " t51_1071 = "& Convert_SLV_To_Hex_String(t51_1071) & " t52_1079 = "& Convert_SLV_To_Hex_String(t52_1079) & " outputs:" & " out5_1087= "  & Convert_SLV_To_Hex_String(out5_1087));
      --
    end process; 
    -- flow-through select operator MUX_1086_inst
    out5_1087 <= t51_1071 when (SGT_i16_u1_1083_wire(0) /=  '0') else t52_1079;
    -- logger for split-operator MUX_1094_inst flow-through 
    process(t61_1095) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1094_inst:flowthrough inputs: " & " SGT_i16_u1_1091_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1091_wire) & " a16_735 = "& Convert_SLV_To_Hex_String(a16_735) & " a26_799 = "& Convert_SLV_To_Hex_String(a26_799) & " outputs:" & " t61_1095= "  & Convert_SLV_To_Hex_String(t61_1095));
      --
    end process; 
    -- flow-through select operator MUX_1094_inst
    t61_1095 <= a16_735 when (SGT_i16_u1_1091_wire(0) /=  '0') else a26_799;
    -- logger for split-operator MUX_1102_inst flow-through 
    process(t62_1103) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1102_inst:flowthrough inputs: " & " SGT_i16_u1_1099_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1099_wire) & " a36_863 = "& Convert_SLV_To_Hex_String(a36_863) & " a46_927 = "& Convert_SLV_To_Hex_String(a46_927) & " outputs:" & " t62_1103= "  & Convert_SLV_To_Hex_String(t62_1103));
      --
    end process; 
    -- flow-through select operator MUX_1102_inst
    t62_1103 <= a36_863 when (SGT_i16_u1_1099_wire(0) /=  '0') else a46_927;
    -- logger for split-operator MUX_1110_inst flow-through 
    process(out6_1111) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1110_inst:flowthrough inputs: " & " SGT_i16_u1_1107_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1107_wire) & " t61_1095 = "& Convert_SLV_To_Hex_String(t61_1095) & " t62_1103 = "& Convert_SLV_To_Hex_String(t62_1103) & " outputs:" & " out6_1111= "  & Convert_SLV_To_Hex_String(out6_1111));
      --
    end process; 
    -- flow-through select operator MUX_1110_inst
    out6_1111 <= t61_1095 when (SGT_i16_u1_1107_wire(0) /=  '0') else t62_1103;
    -- logger for split-operator MUX_1118_inst flow-through 
    process(t71_1119) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1118_inst:flowthrough inputs: " & " SGT_i16_u1_1115_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1115_wire) & " a17_739 = "& Convert_SLV_To_Hex_String(a17_739) & " a27_803 = "& Convert_SLV_To_Hex_String(a27_803) & " outputs:" & " t71_1119= "  & Convert_SLV_To_Hex_String(t71_1119));
      --
    end process; 
    -- flow-through select operator MUX_1118_inst
    t71_1119 <= a17_739 when (SGT_i16_u1_1115_wire(0) /=  '0') else a27_803;
    -- logger for split-operator MUX_1126_inst flow-through 
    process(t72_1127) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1126_inst:flowthrough inputs: " & " SGT_i16_u1_1123_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1123_wire) & " a37_867 = "& Convert_SLV_To_Hex_String(a37_867) & " a47_931 = "& Convert_SLV_To_Hex_String(a47_931) & " outputs:" & " t72_1127= "  & Convert_SLV_To_Hex_String(t72_1127));
      --
    end process; 
    -- flow-through select operator MUX_1126_inst
    t72_1127 <= a37_867 when (SGT_i16_u1_1123_wire(0) /=  '0') else a47_931;
    -- logger for split-operator MUX_1134_inst flow-through 
    process(out7_1135) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1134_inst:flowthrough inputs: " & " SGT_i16_u1_1131_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1131_wire) & " t71_1119 = "& Convert_SLV_To_Hex_String(t71_1119) & " t72_1127 = "& Convert_SLV_To_Hex_String(t72_1127) & " outputs:" & " out7_1135= "  & Convert_SLV_To_Hex_String(out7_1135));
      --
    end process; 
    -- flow-through select operator MUX_1134_inst
    out7_1135 <= t71_1119 when (SGT_i16_u1_1131_wire(0) /=  '0') else t72_1127;
    -- logger for split-operator MUX_1142_inst flow-through 
    process(t81_1143) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1142_inst:flowthrough inputs: " & " SGT_i16_u1_1139_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1139_wire) & " a18_743 = "& Convert_SLV_To_Hex_String(a18_743) & " a28_807 = "& Convert_SLV_To_Hex_String(a28_807) & " outputs:" & " t81_1143= "  & Convert_SLV_To_Hex_String(t81_1143));
      --
    end process; 
    -- flow-through select operator MUX_1142_inst
    t81_1143 <= a18_743 when (SGT_i16_u1_1139_wire(0) /=  '0') else a28_807;
    -- logger for split-operator MUX_1150_inst flow-through 
    process(t82_1151) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1150_inst:flowthrough inputs: " & " SGT_i16_u1_1147_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1147_wire) & " a38_871 = "& Convert_SLV_To_Hex_String(a38_871) & " a48_935 = "& Convert_SLV_To_Hex_String(a48_935) & " outputs:" & " t82_1151= "  & Convert_SLV_To_Hex_String(t82_1151));
      --
    end process; 
    -- flow-through select operator MUX_1150_inst
    t82_1151 <= a38_871 when (SGT_i16_u1_1147_wire(0) /=  '0') else a48_935;
    -- logger for split-operator MUX_1158_inst flow-through 
    process(out8_1159) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1158_inst:flowthrough inputs: " & " SGT_i16_u1_1155_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1155_wire) & " t81_1143 = "& Convert_SLV_To_Hex_String(t81_1143) & " t82_1151 = "& Convert_SLV_To_Hex_String(t82_1151) & " outputs:" & " out8_1159= "  & Convert_SLV_To_Hex_String(out8_1159));
      --
    end process; 
    -- flow-through select operator MUX_1158_inst
    out8_1159 <= t81_1143 when (SGT_i16_u1_1155_wire(0) /=  '0') else t82_1151;
    -- logger for split-operator MUX_1166_inst flow-through 
    process(t91_1167) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1166_inst:flowthrough inputs: " & " SGT_i16_u1_1163_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1163_wire) & " a19_747 = "& Convert_SLV_To_Hex_String(a19_747) & " a29_811 = "& Convert_SLV_To_Hex_String(a29_811) & " outputs:" & " t91_1167= "  & Convert_SLV_To_Hex_String(t91_1167));
      --
    end process; 
    -- flow-through select operator MUX_1166_inst
    t91_1167 <= a19_747 when (SGT_i16_u1_1163_wire(0) /=  '0') else a29_811;
    -- logger for split-operator MUX_1174_inst flow-through 
    process(t92_1175) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1174_inst:flowthrough inputs: " & " SGT_i16_u1_1171_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1171_wire) & " a39_875 = "& Convert_SLV_To_Hex_String(a39_875) & " a49_939 = "& Convert_SLV_To_Hex_String(a49_939) & " outputs:" & " t92_1175= "  & Convert_SLV_To_Hex_String(t92_1175));
      --
    end process; 
    -- flow-through select operator MUX_1174_inst
    t92_1175 <= a39_875 when (SGT_i16_u1_1171_wire(0) /=  '0') else a49_939;
    -- logger for split-operator MUX_1182_inst flow-through 
    process(out9_1183) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1182_inst:flowthrough inputs: " & " SGT_i16_u1_1179_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1179_wire) & " t91_1167 = "& Convert_SLV_To_Hex_String(t91_1167) & " t92_1175 = "& Convert_SLV_To_Hex_String(t92_1175) & " outputs:" & " out9_1183= "  & Convert_SLV_To_Hex_String(out9_1183));
      --
    end process; 
    -- flow-through select operator MUX_1182_inst
    out9_1183 <= t91_1167 when (SGT_i16_u1_1179_wire(0) /=  '0') else t92_1175;
    -- logger for split-operator MUX_1190_inst flow-through 
    process(t101_1191) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1190_inst:flowthrough inputs: " & " SGT_i16_u1_1187_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1187_wire) & " a110_751 = "& Convert_SLV_To_Hex_String(a110_751) & " a210_815 = "& Convert_SLV_To_Hex_String(a210_815) & " outputs:" & " t101_1191= "  & Convert_SLV_To_Hex_String(t101_1191));
      --
    end process; 
    -- flow-through select operator MUX_1190_inst
    t101_1191 <= a110_751 when (SGT_i16_u1_1187_wire(0) /=  '0') else a210_815;
    -- logger for split-operator MUX_1198_inst flow-through 
    process(t102_1199) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1198_inst:flowthrough inputs: " & " SGT_i16_u1_1195_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1195_wire) & " a310_879 = "& Convert_SLV_To_Hex_String(a310_879) & " a410_943 = "& Convert_SLV_To_Hex_String(a410_943) & " outputs:" & " t102_1199= "  & Convert_SLV_To_Hex_String(t102_1199));
      --
    end process; 
    -- flow-through select operator MUX_1198_inst
    t102_1199 <= a310_879 when (SGT_i16_u1_1195_wire(0) /=  '0') else a410_943;
    -- logger for split-operator MUX_1206_inst flow-through 
    process(out10_1207) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1206_inst:flowthrough inputs: " & " SGT_i16_u1_1203_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1203_wire) & " t101_1191 = "& Convert_SLV_To_Hex_String(t101_1191) & " t102_1199 = "& Convert_SLV_To_Hex_String(t102_1199) & " outputs:" & " out10_1207= "  & Convert_SLV_To_Hex_String(out10_1207));
      --
    end process; 
    -- flow-through select operator MUX_1206_inst
    out10_1207 <= t101_1191 when (SGT_i16_u1_1203_wire(0) /=  '0') else t102_1199;
    -- logger for split-operator MUX_1214_inst flow-through 
    process(t111_1215) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1214_inst:flowthrough inputs: " & " SGT_i16_u1_1211_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1211_wire) & " a111_755 = "& Convert_SLV_To_Hex_String(a111_755) & " a211_819 = "& Convert_SLV_To_Hex_String(a211_819) & " outputs:" & " t111_1215= "  & Convert_SLV_To_Hex_String(t111_1215));
      --
    end process; 
    -- flow-through select operator MUX_1214_inst
    t111_1215 <= a111_755 when (SGT_i16_u1_1211_wire(0) /=  '0') else a211_819;
    -- logger for split-operator MUX_1222_inst flow-through 
    process(t112_1223) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1222_inst:flowthrough inputs: " & " SGT_i16_u1_1219_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1219_wire) & " a311_883 = "& Convert_SLV_To_Hex_String(a311_883) & " a411_947 = "& Convert_SLV_To_Hex_String(a411_947) & " outputs:" & " t112_1223= "  & Convert_SLV_To_Hex_String(t112_1223));
      --
    end process; 
    -- flow-through select operator MUX_1222_inst
    t112_1223 <= a311_883 when (SGT_i16_u1_1219_wire(0) /=  '0') else a411_947;
    -- logger for split-operator MUX_1230_inst flow-through 
    process(out11_1231) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1230_inst:flowthrough inputs: " & " SGT_i16_u1_1227_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1227_wire) & " t111_1215 = "& Convert_SLV_To_Hex_String(t111_1215) & " t112_1223 = "& Convert_SLV_To_Hex_String(t112_1223) & " outputs:" & " out11_1231= "  & Convert_SLV_To_Hex_String(out11_1231));
      --
    end process; 
    -- flow-through select operator MUX_1230_inst
    out11_1231 <= t111_1215 when (SGT_i16_u1_1227_wire(0) /=  '0') else t112_1223;
    -- logger for split-operator MUX_1238_inst flow-through 
    process(t121_1239) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1238_inst:flowthrough inputs: " & " SGT_i16_u1_1235_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1235_wire) & " a112_759 = "& Convert_SLV_To_Hex_String(a112_759) & " a212_823 = "& Convert_SLV_To_Hex_String(a212_823) & " outputs:" & " t121_1239= "  & Convert_SLV_To_Hex_String(t121_1239));
      --
    end process; 
    -- flow-through select operator MUX_1238_inst
    t121_1239 <= a112_759 when (SGT_i16_u1_1235_wire(0) /=  '0') else a212_823;
    -- logger for split-operator MUX_1246_inst flow-through 
    process(t122_1247) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1246_inst:flowthrough inputs: " & " SGT_i16_u1_1243_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1243_wire) & " a312_887 = "& Convert_SLV_To_Hex_String(a312_887) & " a412_951 = "& Convert_SLV_To_Hex_String(a412_951) & " outputs:" & " t122_1247= "  & Convert_SLV_To_Hex_String(t122_1247));
      --
    end process; 
    -- flow-through select operator MUX_1246_inst
    t122_1247 <= a312_887 when (SGT_i16_u1_1243_wire(0) /=  '0') else a412_951;
    -- logger for split-operator MUX_1254_inst flow-through 
    process(out12_1255) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1254_inst:flowthrough inputs: " & " SGT_i16_u1_1251_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1251_wire) & " t121_1239 = "& Convert_SLV_To_Hex_String(t121_1239) & " t122_1247 = "& Convert_SLV_To_Hex_String(t122_1247) & " outputs:" & " out12_1255= "  & Convert_SLV_To_Hex_String(out12_1255));
      --
    end process; 
    -- flow-through select operator MUX_1254_inst
    out12_1255 <= t121_1239 when (SGT_i16_u1_1251_wire(0) /=  '0') else t122_1247;
    -- logger for split-operator MUX_1262_inst flow-through 
    process(t131_1263) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1262_inst:flowthrough inputs: " & " SGT_i16_u1_1259_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1259_wire) & " a113_763 = "& Convert_SLV_To_Hex_String(a113_763) & " a213_827 = "& Convert_SLV_To_Hex_String(a213_827) & " outputs:" & " t131_1263= "  & Convert_SLV_To_Hex_String(t131_1263));
      --
    end process; 
    -- flow-through select operator MUX_1262_inst
    t131_1263 <= a113_763 when (SGT_i16_u1_1259_wire(0) /=  '0') else a213_827;
    -- logger for split-operator MUX_1270_inst flow-through 
    process(t132_1271) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1270_inst:flowthrough inputs: " & " SGT_i16_u1_1267_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1267_wire) & " a313_891 = "& Convert_SLV_To_Hex_String(a313_891) & " a413_955 = "& Convert_SLV_To_Hex_String(a413_955) & " outputs:" & " t132_1271= "  & Convert_SLV_To_Hex_String(t132_1271));
      --
    end process; 
    -- flow-through select operator MUX_1270_inst
    t132_1271 <= a313_891 when (SGT_i16_u1_1267_wire(0) /=  '0') else a413_955;
    -- logger for split-operator MUX_1278_inst flow-through 
    process(out13_1279) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1278_inst:flowthrough inputs: " & " SGT_i16_u1_1275_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1275_wire) & " t131_1263 = "& Convert_SLV_To_Hex_String(t131_1263) & " t132_1271 = "& Convert_SLV_To_Hex_String(t132_1271) & " outputs:" & " out13_1279= "  & Convert_SLV_To_Hex_String(out13_1279));
      --
    end process; 
    -- flow-through select operator MUX_1278_inst
    out13_1279 <= t131_1263 when (SGT_i16_u1_1275_wire(0) /=  '0') else t132_1271;
    -- logger for split-operator MUX_1286_inst flow-through 
    process(t141_1287) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1286_inst:flowthrough inputs: " & " SGT_i16_u1_1283_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1283_wire) & " a114_767 = "& Convert_SLV_To_Hex_String(a114_767) & " a214_831 = "& Convert_SLV_To_Hex_String(a214_831) & " outputs:" & " t141_1287= "  & Convert_SLV_To_Hex_String(t141_1287));
      --
    end process; 
    -- flow-through select operator MUX_1286_inst
    t141_1287 <= a114_767 when (SGT_i16_u1_1283_wire(0) /=  '0') else a214_831;
    -- logger for split-operator MUX_1294_inst flow-through 
    process(t142_1295) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1294_inst:flowthrough inputs: " & " SGT_i16_u1_1291_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1291_wire) & " a314_895 = "& Convert_SLV_To_Hex_String(a314_895) & " a414_959 = "& Convert_SLV_To_Hex_String(a414_959) & " outputs:" & " t142_1295= "  & Convert_SLV_To_Hex_String(t142_1295));
      --
    end process; 
    -- flow-through select operator MUX_1294_inst
    t142_1295 <= a314_895 when (SGT_i16_u1_1291_wire(0) /=  '0') else a414_959;
    -- logger for split-operator MUX_1302_inst flow-through 
    process(out14_1303) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1302_inst:flowthrough inputs: " & " SGT_i16_u1_1299_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1299_wire) & " t141_1287 = "& Convert_SLV_To_Hex_String(t141_1287) & " t142_1295 = "& Convert_SLV_To_Hex_String(t142_1295) & " outputs:" & " out14_1303= "  & Convert_SLV_To_Hex_String(out14_1303));
      --
    end process; 
    -- flow-through select operator MUX_1302_inst
    out14_1303 <= t141_1287 when (SGT_i16_u1_1299_wire(0) /=  '0') else t142_1295;
    -- logger for split-operator MUX_1310_inst flow-through 
    process(t151_1311) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1310_inst:flowthrough inputs: " & " SGT_i16_u1_1307_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1307_wire) & " a115_771 = "& Convert_SLV_To_Hex_String(a115_771) & " a215_835 = "& Convert_SLV_To_Hex_String(a215_835) & " outputs:" & " t151_1311= "  & Convert_SLV_To_Hex_String(t151_1311));
      --
    end process; 
    -- flow-through select operator MUX_1310_inst
    t151_1311 <= a115_771 when (SGT_i16_u1_1307_wire(0) /=  '0') else a215_835;
    -- logger for split-operator MUX_1318_inst flow-through 
    process(t152_1319) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1318_inst:flowthrough inputs: " & " SGT_i16_u1_1315_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1315_wire) & " a315_899 = "& Convert_SLV_To_Hex_String(a315_899) & " a415_963 = "& Convert_SLV_To_Hex_String(a415_963) & " outputs:" & " t152_1319= "  & Convert_SLV_To_Hex_String(t152_1319));
      --
    end process; 
    -- flow-through select operator MUX_1318_inst
    t152_1319 <= a315_899 when (SGT_i16_u1_1315_wire(0) /=  '0') else a415_963;
    -- logger for split-operator MUX_1326_inst flow-through 
    process(out15_1327) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1326_inst:flowthrough inputs: " & " SGT_i16_u1_1323_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1323_wire) & " t151_1311 = "& Convert_SLV_To_Hex_String(t151_1311) & " t152_1319 = "& Convert_SLV_To_Hex_String(t152_1319) & " outputs:" & " out15_1327= "  & Convert_SLV_To_Hex_String(out15_1327));
      --
    end process; 
    -- flow-through select operator MUX_1326_inst
    out15_1327 <= t151_1311 when (SGT_i16_u1_1323_wire(0) /=  '0') else t152_1319;
    -- logger for split-operator MUX_1334_inst flow-through 
    process(t161_1335) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1334_inst:flowthrough inputs: " & " SGT_i16_u1_1331_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1331_wire) & " a116_775 = "& Convert_SLV_To_Hex_String(a116_775) & " a216_839 = "& Convert_SLV_To_Hex_String(a216_839) & " outputs:" & " t161_1335= "  & Convert_SLV_To_Hex_String(t161_1335));
      --
    end process; 
    -- flow-through select operator MUX_1334_inst
    t161_1335 <= a116_775 when (SGT_i16_u1_1331_wire(0) /=  '0') else a216_839;
    -- logger for split-operator MUX_1342_inst flow-through 
    process(t162_1343) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1342_inst:flowthrough inputs: " & " SGT_i16_u1_1339_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1339_wire) & " a316_903 = "& Convert_SLV_To_Hex_String(a316_903) & " a416_967 = "& Convert_SLV_To_Hex_String(a416_967) & " outputs:" & " t162_1343= "  & Convert_SLV_To_Hex_String(t162_1343));
      --
    end process; 
    -- flow-through select operator MUX_1342_inst
    t162_1343 <= a316_903 when (SGT_i16_u1_1339_wire(0) /=  '0') else a416_967;
    -- logger for split-operator MUX_1350_inst flow-through 
    process(out16_1351) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_1350_inst:flowthrough inputs: " & " SGT_i16_u1_1347_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_1347_wire) & " t161_1335 = "& Convert_SLV_To_Hex_String(t161_1335) & " t162_1343 = "& Convert_SLV_To_Hex_String(t162_1343) & " outputs:" & " out16_1351= "  & Convert_SLV_To_Hex_String(out16_1351));
      --
    end process; 
    -- flow-through select operator MUX_1350_inst
    out16_1351 <= t161_1335 when (SGT_i16_u1_1347_wire(0) /=  '0') else t162_1343;
    -- logger for split-operator MUX_974_inst flow-through 
    process(t11_975) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_974_inst:flowthrough inputs: " & " SGT_i16_u1_971_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_971_wire) & " a11_715 = "& Convert_SLV_To_Hex_String(a11_715) & " a21_779 = "& Convert_SLV_To_Hex_String(a21_779) & " outputs:" & " t11_975= "  & Convert_SLV_To_Hex_String(t11_975));
      --
    end process; 
    -- flow-through select operator MUX_974_inst
    t11_975 <= a11_715 when (SGT_i16_u1_971_wire(0) /=  '0') else a21_779;
    -- logger for split-operator MUX_982_inst flow-through 
    process(t12_983) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_982_inst:flowthrough inputs: " & " SGT_i16_u1_979_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_979_wire) & " a31_843 = "& Convert_SLV_To_Hex_String(a31_843) & " a41_907 = "& Convert_SLV_To_Hex_String(a41_907) & " outputs:" & " t12_983= "  & Convert_SLV_To_Hex_String(t12_983));
      --
    end process; 
    -- flow-through select operator MUX_982_inst
    t12_983 <= a31_843 when (SGT_i16_u1_979_wire(0) /=  '0') else a41_907;
    -- logger for split-operator MUX_990_inst flow-through 
    process(out1_991) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_990_inst:flowthrough inputs: " & " SGT_i16_u1_987_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_987_wire) & " t11_975 = "& Convert_SLV_To_Hex_String(t11_975) & " t12_983 = "& Convert_SLV_To_Hex_String(t12_983) & " outputs:" & " out1_991= "  & Convert_SLV_To_Hex_String(out1_991));
      --
    end process; 
    -- flow-through select operator MUX_990_inst
    out1_991 <= t11_975 when (SGT_i16_u1_987_wire(0) /=  '0') else t12_983;
    -- logger for split-operator MUX_998_inst flow-through 
    process(t21_999) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:MUX_998_inst:flowthrough inputs: " & " SGT_i16_u1_995_wire = "& Convert_SLV_To_Hex_String(SGT_i16_u1_995_wire) & " a12_719 = "& Convert_SLV_To_Hex_String(a12_719) & " a22_783 = "& Convert_SLV_To_Hex_String(a22_783) & " outputs:" & " t21_999= "  & Convert_SLV_To_Hex_String(t21_999));
      --
    end process; 
    -- flow-through select operator MUX_998_inst
    t21_999 <= a12_719 when (SGT_i16_u1_995_wire(0) /=  '0') else a22_783;
    -- logger for split-operator slice_457_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_457_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_457_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_457_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_457_inst:finished:  outputs: " & " sliced_v11_458= "  & Convert_SLV_To_Hex_String(sliced_v11_458));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_457_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_457_inst_req_0;
      slice_457_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_457_inst_req_1;
      slice_457_inst_ack_1<= update_ack(0);
      slice_457_inst: SliceSplitProtocol generic map(name => "slice_457_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v11_458, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_461_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_461_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_461_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_461_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_461_inst:finished:  outputs: " & " sliced_v12_462= "  & Convert_SLV_To_Hex_String(sliced_v12_462));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_461_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_461_inst_req_0;
      slice_461_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_461_inst_req_1;
      slice_461_inst_ack_1<= update_ack(0);
      slice_461_inst: SliceSplitProtocol generic map(name => "slice_461_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v12_462, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_465_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_465_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_465_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_465_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_465_inst:finished:  outputs: " & " sliced_v13_466= "  & Convert_SLV_To_Hex_String(sliced_v13_466));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_465_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_465_inst_req_0;
      slice_465_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_465_inst_req_1;
      slice_465_inst_ack_1<= update_ack(0);
      slice_465_inst: SliceSplitProtocol generic map(name => "slice_465_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v13_466, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_469_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_469_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_469_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_469_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_469_inst:finished:  outputs: " & " sliced_v14_470= "  & Convert_SLV_To_Hex_String(sliced_v14_470));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_469_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_469_inst_req_0;
      slice_469_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_469_inst_req_1;
      slice_469_inst_ack_1<= update_ack(0);
      slice_469_inst: SliceSplitProtocol generic map(name => "slice_469_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v14_470, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_473_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_473_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_473_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_473_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_473_inst:finished:  outputs: " & " sliced_v15_474= "  & Convert_SLV_To_Hex_String(sliced_v15_474));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_473_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_473_inst_req_0;
      slice_473_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_473_inst_req_1;
      slice_473_inst_ack_1<= update_ack(0);
      slice_473_inst: SliceSplitProtocol generic map(name => "slice_473_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v15_474, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_477_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_477_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_477_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_477_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_477_inst:finished:  outputs: " & " sliced_v16_478= "  & Convert_SLV_To_Hex_String(sliced_v16_478));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_477_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_477_inst_req_0;
      slice_477_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_477_inst_req_1;
      slice_477_inst_ack_1<= update_ack(0);
      slice_477_inst: SliceSplitProtocol generic map(name => "slice_477_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v16_478, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_481_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_481_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_481_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_481_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_481_inst:finished:  outputs: " & " sliced_v17_482= "  & Convert_SLV_To_Hex_String(sliced_v17_482));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_481_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_481_inst_req_0;
      slice_481_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_481_inst_req_1;
      slice_481_inst_ack_1<= update_ack(0);
      slice_481_inst: SliceSplitProtocol generic map(name => "slice_481_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v17_482, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_485_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_485_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_485_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_485_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_485_inst:finished:  outputs: " & " sliced_v18_486= "  & Convert_SLV_To_Hex_String(sliced_v18_486));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_485_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_485_inst_req_0;
      slice_485_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_485_inst_req_1;
      slice_485_inst_ack_1<= update_ack(0);
      slice_485_inst: SliceSplitProtocol generic map(name => "slice_485_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v18_486, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_489_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_489_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_489_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_489_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_489_inst:finished:  outputs: " & " sliced_v19_490= "  & Convert_SLV_To_Hex_String(sliced_v19_490));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_489_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_489_inst_req_0;
      slice_489_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_489_inst_req_1;
      slice_489_inst_ack_1<= update_ack(0);
      slice_489_inst: SliceSplitProtocol generic map(name => "slice_489_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v19_490, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_493_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_493_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_493_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_493_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_493_inst:finished:  outputs: " & " sliced_v110_494= "  & Convert_SLV_To_Hex_String(sliced_v110_494));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_493_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_493_inst_req_0;
      slice_493_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_493_inst_req_1;
      slice_493_inst_ack_1<= update_ack(0);
      slice_493_inst: SliceSplitProtocol generic map(name => "slice_493_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v110_494, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_497_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_497_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_497_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_497_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_497_inst:finished:  outputs: " & " sliced_v111_498= "  & Convert_SLV_To_Hex_String(sliced_v111_498));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_497_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_497_inst_req_0;
      slice_497_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_497_inst_req_1;
      slice_497_inst_ack_1<= update_ack(0);
      slice_497_inst: SliceSplitProtocol generic map(name => "slice_497_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v111_498, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_501_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_501_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_501_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_501_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_501_inst:finished:  outputs: " & " sliced_v112_502= "  & Convert_SLV_To_Hex_String(sliced_v112_502));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_501_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_501_inst_req_0;
      slice_501_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_501_inst_req_1;
      slice_501_inst_ack_1<= update_ack(0);
      slice_501_inst: SliceSplitProtocol generic map(name => "slice_501_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v112_502, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_505_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_505_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_505_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_505_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_505_inst:finished:  outputs: " & " sliced_v113_506= "  & Convert_SLV_To_Hex_String(sliced_v113_506));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_505_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_505_inst_req_0;
      slice_505_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_505_inst_req_1;
      slice_505_inst_ack_1<= update_ack(0);
      slice_505_inst: SliceSplitProtocol generic map(name => "slice_505_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v113_506, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_509_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_509_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_509_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_509_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_509_inst:finished:  outputs: " & " sliced_v114_510= "  & Convert_SLV_To_Hex_String(sliced_v114_510));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_509_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_509_inst_req_0;
      slice_509_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_509_inst_req_1;
      slice_509_inst_ack_1<= update_ack(0);
      slice_509_inst: SliceSplitProtocol generic map(name => "slice_509_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v114_510, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_513_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_513_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_513_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_513_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_513_inst:finished:  outputs: " & " sliced_v115_514= "  & Convert_SLV_To_Hex_String(sliced_v115_514));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_513_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_513_inst_req_0;
      slice_513_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_513_inst_req_1;
      slice_513_inst_ack_1<= update_ack(0);
      slice_513_inst: SliceSplitProtocol generic map(name => "slice_513_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v115_514, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_517_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_517_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_517_inst:started:   inputs: " & " c1_442 = "& Convert_SLV_To_Hex_String(c1_442));
          --
        end if; 
        if slice_517_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_517_inst:finished:  outputs: " & " sliced_v116_518= "  & Convert_SLV_To_Hex_String(sliced_v116_518));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_517_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_517_inst_req_0;
      slice_517_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_517_inst_req_1;
      slice_517_inst_ack_1<= update_ack(0);
      slice_517_inst: SliceSplitProtocol generic map(name => "slice_517_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_442, dout => sliced_v116_518, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_521_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_521_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_521_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_521_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_521_inst:finished:  outputs: " & " sliced_v21_522= "  & Convert_SLV_To_Hex_String(sliced_v21_522));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_521_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_521_inst_req_0;
      slice_521_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_521_inst_req_1;
      slice_521_inst_ack_1<= update_ack(0);
      slice_521_inst: SliceSplitProtocol generic map(name => "slice_521_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v21_522, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_525_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_525_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_525_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_525_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_525_inst:finished:  outputs: " & " sliced_v22_526= "  & Convert_SLV_To_Hex_String(sliced_v22_526));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_525_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_525_inst_req_0;
      slice_525_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_525_inst_req_1;
      slice_525_inst_ack_1<= update_ack(0);
      slice_525_inst: SliceSplitProtocol generic map(name => "slice_525_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v22_526, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_529_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_529_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_529_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_529_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_529_inst:finished:  outputs: " & " sliced_v23_530= "  & Convert_SLV_To_Hex_String(sliced_v23_530));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_529_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_529_inst_req_0;
      slice_529_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_529_inst_req_1;
      slice_529_inst_ack_1<= update_ack(0);
      slice_529_inst: SliceSplitProtocol generic map(name => "slice_529_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v23_530, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_533_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_533_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_533_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_533_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_533_inst:finished:  outputs: " & " sliced_v24_534= "  & Convert_SLV_To_Hex_String(sliced_v24_534));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_533_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_533_inst_req_0;
      slice_533_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_533_inst_req_1;
      slice_533_inst_ack_1<= update_ack(0);
      slice_533_inst: SliceSplitProtocol generic map(name => "slice_533_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v24_534, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_537_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_537_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_537_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_537_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_537_inst:finished:  outputs: " & " sliced_v25_538= "  & Convert_SLV_To_Hex_String(sliced_v25_538));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_537_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_537_inst_req_0;
      slice_537_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_537_inst_req_1;
      slice_537_inst_ack_1<= update_ack(0);
      slice_537_inst: SliceSplitProtocol generic map(name => "slice_537_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v25_538, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_541_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_541_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_541_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_541_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_541_inst:finished:  outputs: " & " sliced_v26_542= "  & Convert_SLV_To_Hex_String(sliced_v26_542));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_541_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_541_inst_req_0;
      slice_541_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_541_inst_req_1;
      slice_541_inst_ack_1<= update_ack(0);
      slice_541_inst: SliceSplitProtocol generic map(name => "slice_541_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v26_542, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_545_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_545_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_545_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_545_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_545_inst:finished:  outputs: " & " sliced_v27_546= "  & Convert_SLV_To_Hex_String(sliced_v27_546));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_545_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_545_inst_req_0;
      slice_545_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_545_inst_req_1;
      slice_545_inst_ack_1<= update_ack(0);
      slice_545_inst: SliceSplitProtocol generic map(name => "slice_545_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v27_546, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_549_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_549_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_549_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_549_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_549_inst:finished:  outputs: " & " sliced_v28_550= "  & Convert_SLV_To_Hex_String(sliced_v28_550));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_549_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_549_inst_req_0;
      slice_549_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_549_inst_req_1;
      slice_549_inst_ack_1<= update_ack(0);
      slice_549_inst: SliceSplitProtocol generic map(name => "slice_549_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v28_550, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_553_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_553_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_553_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_553_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_553_inst:finished:  outputs: " & " sliced_v29_554= "  & Convert_SLV_To_Hex_String(sliced_v29_554));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_553_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_553_inst_req_0;
      slice_553_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_553_inst_req_1;
      slice_553_inst_ack_1<= update_ack(0);
      slice_553_inst: SliceSplitProtocol generic map(name => "slice_553_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v29_554, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_557_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_557_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_557_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_557_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_557_inst:finished:  outputs: " & " sliced_v210_558= "  & Convert_SLV_To_Hex_String(sliced_v210_558));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_557_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_557_inst_req_0;
      slice_557_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_557_inst_req_1;
      slice_557_inst_ack_1<= update_ack(0);
      slice_557_inst: SliceSplitProtocol generic map(name => "slice_557_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v210_558, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_561_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_561_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_561_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_561_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_561_inst:finished:  outputs: " & " sliced_v211_562= "  & Convert_SLV_To_Hex_String(sliced_v211_562));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_561_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_561_inst_req_0;
      slice_561_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_561_inst_req_1;
      slice_561_inst_ack_1<= update_ack(0);
      slice_561_inst: SliceSplitProtocol generic map(name => "slice_561_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v211_562, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_565_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_565_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_565_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_565_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_565_inst:finished:  outputs: " & " sliced_v212_566= "  & Convert_SLV_To_Hex_String(sliced_v212_566));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_565_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_565_inst_req_0;
      slice_565_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_565_inst_req_1;
      slice_565_inst_ack_1<= update_ack(0);
      slice_565_inst: SliceSplitProtocol generic map(name => "slice_565_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v212_566, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_569_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_569_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_569_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_569_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_569_inst:finished:  outputs: " & " sliced_v213_570= "  & Convert_SLV_To_Hex_String(sliced_v213_570));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_569_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_569_inst_req_0;
      slice_569_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_569_inst_req_1;
      slice_569_inst_ack_1<= update_ack(0);
      slice_569_inst: SliceSplitProtocol generic map(name => "slice_569_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v213_570, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_573_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_573_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_573_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_573_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_573_inst:finished:  outputs: " & " sliced_v214_574= "  & Convert_SLV_To_Hex_String(sliced_v214_574));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_573_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_573_inst_req_0;
      slice_573_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_573_inst_req_1;
      slice_573_inst_ack_1<= update_ack(0);
      slice_573_inst: SliceSplitProtocol generic map(name => "slice_573_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v214_574, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_577_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_577_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_577_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_577_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_577_inst:finished:  outputs: " & " sliced_v215_578= "  & Convert_SLV_To_Hex_String(sliced_v215_578));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_577_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_577_inst_req_0;
      slice_577_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_577_inst_req_1;
      slice_577_inst_ack_1<= update_ack(0);
      slice_577_inst: SliceSplitProtocol generic map(name => "slice_577_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v215_578, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_581_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_581_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_581_inst:started:   inputs: " & " c2_446 = "& Convert_SLV_To_Hex_String(c2_446));
          --
        end if; 
        if slice_581_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_581_inst:finished:  outputs: " & " sliced_v216_582= "  & Convert_SLV_To_Hex_String(sliced_v216_582));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_581_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_581_inst_req_0;
      slice_581_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_581_inst_req_1;
      slice_581_inst_ack_1<= update_ack(0);
      slice_581_inst: SliceSplitProtocol generic map(name => "slice_581_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_446, dout => sliced_v216_582, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_585_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_585_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_585_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_585_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_585_inst:finished:  outputs: " & " sliced_v31_586= "  & Convert_SLV_To_Hex_String(sliced_v31_586));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_585_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_585_inst_req_0;
      slice_585_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_585_inst_req_1;
      slice_585_inst_ack_1<= update_ack(0);
      slice_585_inst: SliceSplitProtocol generic map(name => "slice_585_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v31_586, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_589_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_589_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_589_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_589_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_589_inst:finished:  outputs: " & " sliced_v32_590= "  & Convert_SLV_To_Hex_String(sliced_v32_590));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_589_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_589_inst_req_0;
      slice_589_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_589_inst_req_1;
      slice_589_inst_ack_1<= update_ack(0);
      slice_589_inst: SliceSplitProtocol generic map(name => "slice_589_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v32_590, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_593_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_593_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_593_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_593_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_593_inst:finished:  outputs: " & " sliced_v33_594= "  & Convert_SLV_To_Hex_String(sliced_v33_594));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_593_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_593_inst_req_0;
      slice_593_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_593_inst_req_1;
      slice_593_inst_ack_1<= update_ack(0);
      slice_593_inst: SliceSplitProtocol generic map(name => "slice_593_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v33_594, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_597_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_597_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_597_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_597_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_597_inst:finished:  outputs: " & " sliced_v34_598= "  & Convert_SLV_To_Hex_String(sliced_v34_598));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_597_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_597_inst_req_0;
      slice_597_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_597_inst_req_1;
      slice_597_inst_ack_1<= update_ack(0);
      slice_597_inst: SliceSplitProtocol generic map(name => "slice_597_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v34_598, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_601_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_601_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_601_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_601_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_601_inst:finished:  outputs: " & " sliced_v35_602= "  & Convert_SLV_To_Hex_String(sliced_v35_602));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_601_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_601_inst_req_0;
      slice_601_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_601_inst_req_1;
      slice_601_inst_ack_1<= update_ack(0);
      slice_601_inst: SliceSplitProtocol generic map(name => "slice_601_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v35_602, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_605_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_605_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_605_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_605_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_605_inst:finished:  outputs: " & " sliced_v36_606= "  & Convert_SLV_To_Hex_String(sliced_v36_606));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_605_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_605_inst_req_0;
      slice_605_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_605_inst_req_1;
      slice_605_inst_ack_1<= update_ack(0);
      slice_605_inst: SliceSplitProtocol generic map(name => "slice_605_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v36_606, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_609_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_609_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_609_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_609_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_609_inst:finished:  outputs: " & " sliced_v37_610= "  & Convert_SLV_To_Hex_String(sliced_v37_610));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_609_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_609_inst_req_0;
      slice_609_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_609_inst_req_1;
      slice_609_inst_ack_1<= update_ack(0);
      slice_609_inst: SliceSplitProtocol generic map(name => "slice_609_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v37_610, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_613_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_613_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_613_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_613_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_613_inst:finished:  outputs: " & " sliced_v38_614= "  & Convert_SLV_To_Hex_String(sliced_v38_614));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_613_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_613_inst_req_0;
      slice_613_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_613_inst_req_1;
      slice_613_inst_ack_1<= update_ack(0);
      slice_613_inst: SliceSplitProtocol generic map(name => "slice_613_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v38_614, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_617_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_617_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_617_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_617_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_617_inst:finished:  outputs: " & " sliced_v39_618= "  & Convert_SLV_To_Hex_String(sliced_v39_618));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_617_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_617_inst_req_0;
      slice_617_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_617_inst_req_1;
      slice_617_inst_ack_1<= update_ack(0);
      slice_617_inst: SliceSplitProtocol generic map(name => "slice_617_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v39_618, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_621_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_621_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_621_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_621_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_621_inst:finished:  outputs: " & " sliced_v310_622= "  & Convert_SLV_To_Hex_String(sliced_v310_622));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_621_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_621_inst_req_0;
      slice_621_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_621_inst_req_1;
      slice_621_inst_ack_1<= update_ack(0);
      slice_621_inst: SliceSplitProtocol generic map(name => "slice_621_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v310_622, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_625_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_625_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_625_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_625_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_625_inst:finished:  outputs: " & " sliced_v311_626= "  & Convert_SLV_To_Hex_String(sliced_v311_626));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_625_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_625_inst_req_0;
      slice_625_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_625_inst_req_1;
      slice_625_inst_ack_1<= update_ack(0);
      slice_625_inst: SliceSplitProtocol generic map(name => "slice_625_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v311_626, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_629_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_629_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_629_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_629_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_629_inst:finished:  outputs: " & " sliced_v312_630= "  & Convert_SLV_To_Hex_String(sliced_v312_630));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_629_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_629_inst_req_0;
      slice_629_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_629_inst_req_1;
      slice_629_inst_ack_1<= update_ack(0);
      slice_629_inst: SliceSplitProtocol generic map(name => "slice_629_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v312_630, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_633_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_633_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_633_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_633_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_633_inst:finished:  outputs: " & " sliced_v313_634= "  & Convert_SLV_To_Hex_String(sliced_v313_634));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_633_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_633_inst_req_0;
      slice_633_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_633_inst_req_1;
      slice_633_inst_ack_1<= update_ack(0);
      slice_633_inst: SliceSplitProtocol generic map(name => "slice_633_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v313_634, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_637_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_637_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_637_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_637_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_637_inst:finished:  outputs: " & " sliced_v314_638= "  & Convert_SLV_To_Hex_String(sliced_v314_638));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_637_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_637_inst_req_0;
      slice_637_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_637_inst_req_1;
      slice_637_inst_ack_1<= update_ack(0);
      slice_637_inst: SliceSplitProtocol generic map(name => "slice_637_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v314_638, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_641_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_641_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_641_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_641_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_641_inst:finished:  outputs: " & " sliced_v315_642= "  & Convert_SLV_To_Hex_String(sliced_v315_642));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_641_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_641_inst_req_0;
      slice_641_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_641_inst_req_1;
      slice_641_inst_ack_1<= update_ack(0);
      slice_641_inst: SliceSplitProtocol generic map(name => "slice_641_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v315_642, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_645_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_645_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_645_inst:started:   inputs: " & " c3_450 = "& Convert_SLV_To_Hex_String(c3_450));
          --
        end if; 
        if slice_645_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_645_inst:finished:  outputs: " & " sliced_v316_646= "  & Convert_SLV_To_Hex_String(sliced_v316_646));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_645_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_645_inst_req_0;
      slice_645_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_645_inst_req_1;
      slice_645_inst_ack_1<= update_ack(0);
      slice_645_inst: SliceSplitProtocol generic map(name => "slice_645_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_450, dout => sliced_v316_646, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_649_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_649_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_649_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_649_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_649_inst:finished:  outputs: " & " sliced_v41_650= "  & Convert_SLV_To_Hex_String(sliced_v41_650));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_649_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_649_inst_req_0;
      slice_649_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_649_inst_req_1;
      slice_649_inst_ack_1<= update_ack(0);
      slice_649_inst: SliceSplitProtocol generic map(name => "slice_649_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v41_650, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_653_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_653_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_653_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_653_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_653_inst:finished:  outputs: " & " sliced_v42_654= "  & Convert_SLV_To_Hex_String(sliced_v42_654));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_653_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_653_inst_req_0;
      slice_653_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_653_inst_req_1;
      slice_653_inst_ack_1<= update_ack(0);
      slice_653_inst: SliceSplitProtocol generic map(name => "slice_653_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v42_654, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_657_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_657_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_657_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_657_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_657_inst:finished:  outputs: " & " sliced_v43_658= "  & Convert_SLV_To_Hex_String(sliced_v43_658));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_657_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_657_inst_req_0;
      slice_657_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_657_inst_req_1;
      slice_657_inst_ack_1<= update_ack(0);
      slice_657_inst: SliceSplitProtocol generic map(name => "slice_657_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v43_658, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_661_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_661_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_661_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_661_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_661_inst:finished:  outputs: " & " sliced_v44_662= "  & Convert_SLV_To_Hex_String(sliced_v44_662));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_661_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_661_inst_req_0;
      slice_661_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_661_inst_req_1;
      slice_661_inst_ack_1<= update_ack(0);
      slice_661_inst: SliceSplitProtocol generic map(name => "slice_661_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v44_662, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_665_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_665_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_665_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_665_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_665_inst:finished:  outputs: " & " sliced_v45_666= "  & Convert_SLV_To_Hex_String(sliced_v45_666));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_665_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_665_inst_req_0;
      slice_665_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_665_inst_req_1;
      slice_665_inst_ack_1<= update_ack(0);
      slice_665_inst: SliceSplitProtocol generic map(name => "slice_665_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v45_666, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_669_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_669_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_669_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_669_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_669_inst:finished:  outputs: " & " sliced_v46_670= "  & Convert_SLV_To_Hex_String(sliced_v46_670));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_669_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_669_inst_req_0;
      slice_669_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_669_inst_req_1;
      slice_669_inst_ack_1<= update_ack(0);
      slice_669_inst: SliceSplitProtocol generic map(name => "slice_669_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v46_670, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_673_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_673_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_673_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_673_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_673_inst:finished:  outputs: " & " sliced_v47_674= "  & Convert_SLV_To_Hex_String(sliced_v47_674));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_673_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_673_inst_req_0;
      slice_673_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_673_inst_req_1;
      slice_673_inst_ack_1<= update_ack(0);
      slice_673_inst: SliceSplitProtocol generic map(name => "slice_673_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v47_674, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_677_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_677_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_677_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_677_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_677_inst:finished:  outputs: " & " sliced_v48_678= "  & Convert_SLV_To_Hex_String(sliced_v48_678));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_677_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_677_inst_req_0;
      slice_677_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_677_inst_req_1;
      slice_677_inst_ack_1<= update_ack(0);
      slice_677_inst: SliceSplitProtocol generic map(name => "slice_677_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v48_678, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_681_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_681_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_681_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_681_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_681_inst:finished:  outputs: " & " sliced_v49_682= "  & Convert_SLV_To_Hex_String(sliced_v49_682));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_681_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_681_inst_req_0;
      slice_681_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_681_inst_req_1;
      slice_681_inst_ack_1<= update_ack(0);
      slice_681_inst: SliceSplitProtocol generic map(name => "slice_681_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v49_682, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_685_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_685_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_685_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_685_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_685_inst:finished:  outputs: " & " sliced_v410_686= "  & Convert_SLV_To_Hex_String(sliced_v410_686));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_685_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_685_inst_req_0;
      slice_685_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_685_inst_req_1;
      slice_685_inst_ack_1<= update_ack(0);
      slice_685_inst: SliceSplitProtocol generic map(name => "slice_685_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v410_686, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_689_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_689_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_689_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_689_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_689_inst:finished:  outputs: " & " sliced_v411_690= "  & Convert_SLV_To_Hex_String(sliced_v411_690));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_689_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_689_inst_req_0;
      slice_689_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_689_inst_req_1;
      slice_689_inst_ack_1<= update_ack(0);
      slice_689_inst: SliceSplitProtocol generic map(name => "slice_689_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v411_690, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_693_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_693_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_693_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_693_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_693_inst:finished:  outputs: " & " sliced_v412_694= "  & Convert_SLV_To_Hex_String(sliced_v412_694));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_693_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_693_inst_req_0;
      slice_693_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_693_inst_req_1;
      slice_693_inst_ack_1<= update_ack(0);
      slice_693_inst: SliceSplitProtocol generic map(name => "slice_693_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v412_694, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_697_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_697_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_697_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_697_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_697_inst:finished:  outputs: " & " sliced_v413_698= "  & Convert_SLV_To_Hex_String(sliced_v413_698));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_697_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_697_inst_req_0;
      slice_697_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_697_inst_req_1;
      slice_697_inst_ack_1<= update_ack(0);
      slice_697_inst: SliceSplitProtocol generic map(name => "slice_697_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v413_698, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_701_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_701_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_701_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_701_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_701_inst:finished:  outputs: " & " sliced_v414_702= "  & Convert_SLV_To_Hex_String(sliced_v414_702));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_701_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_701_inst_req_0;
      slice_701_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_701_inst_req_1;
      slice_701_inst_ack_1<= update_ack(0);
      slice_701_inst: SliceSplitProtocol generic map(name => "slice_701_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v414_702, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_705_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_705_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_705_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_705_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_705_inst:finished:  outputs: " & " sliced_v415_706= "  & Convert_SLV_To_Hex_String(sliced_v415_706));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_705_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_705_inst_req_0;
      slice_705_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_705_inst_req_1;
      slice_705_inst_ack_1<= update_ack(0);
      slice_705_inst: SliceSplitProtocol generic map(name => "slice_705_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v415_706, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_709_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_709_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_709_inst:started:   inputs: " & " c4_454 = "& Convert_SLV_To_Hex_String(c4_454));
          --
        end if; 
        if slice_709_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:slice_709_inst:finished:  outputs: " & " sliced_v416_710= "  & Convert_SLV_To_Hex_String(sliced_v416_710));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_709_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_709_inst_req_0;
      slice_709_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_709_inst_req_1;
      slice_709_inst_ack_1<= update_ack(0);
      slice_709_inst: SliceSplitProtocol generic map(name => "slice_709_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_454, dout => sliced_v416_710, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator W_myptr5_1359_delayed_8_0_1359_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_myptr5_1359_delayed_8_0_1359_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:W_myptr5_1359_delayed_8_0_1359_inst:started:   inputs: " & " myptr5_1358 = "& Convert_SLV_To_Hex_String(myptr5_1358));
          --
        end if; 
        if W_myptr5_1359_delayed_8_0_1359_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:W_myptr5_1359_delayed_8_0_1359_inst:finished:  outputs: " & " myptr5_1359_delayed_8_0_1361= "  & Convert_SLV_To_Hex_String(myptr5_1359_delayed_8_0_1361));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_myptr5_1359_delayed_8_0_1359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr5_1359_delayed_8_0_1359_inst_req_0;
      W_myptr5_1359_delayed_8_0_1359_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr5_1359_delayed_8_0_1359_inst_req_1;
      W_myptr5_1359_delayed_8_0_1359_inst_ack_1<= rack(0);
      W_myptr5_1359_delayed_8_0_1359_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr5_1359_delayed_8_0_1359_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr5_1358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr5_1359_delayed_8_0_1361,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_myptr6_1382_delayed_8_0_1385_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_myptr6_1382_delayed_8_0_1385_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:W_myptr6_1382_delayed_8_0_1385_inst:started:   inputs: " & " myptr6_1384 = "& Convert_SLV_To_Hex_String(myptr6_1384));
          --
        end if; 
        if W_myptr6_1382_delayed_8_0_1385_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:W_myptr6_1382_delayed_8_0_1385_inst:finished:  outputs: " & " myptr6_1382_delayed_8_0_1387= "  & Convert_SLV_To_Hex_String(myptr6_1382_delayed_8_0_1387));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_myptr6_1382_delayed_8_0_1385_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr6_1382_delayed_8_0_1385_inst_req_0;
      W_myptr6_1382_delayed_8_0_1385_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr6_1382_delayed_8_0_1385_inst_req_1;
      W_myptr6_1382_delayed_8_0_1385_inst_ack_1<= rack(0);
      W_myptr6_1382_delayed_8_0_1385_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr6_1382_delayed_8_0_1385_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr6_1384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr6_1382_delayed_8_0_1387,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_myptr7_1405_delayed_8_0_1411_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_myptr7_1405_delayed_8_0_1411_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:W_myptr7_1405_delayed_8_0_1411_inst:started:   inputs: " & " myptr7_1410 = "& Convert_SLV_To_Hex_String(myptr7_1410));
          --
        end if; 
        if W_myptr7_1405_delayed_8_0_1411_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:W_myptr7_1405_delayed_8_0_1411_inst:finished:  outputs: " & " myptr7_1405_delayed_8_0_1413= "  & Convert_SLV_To_Hex_String(myptr7_1405_delayed_8_0_1413));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_myptr7_1405_delayed_8_0_1411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr7_1405_delayed_8_0_1411_inst_req_0;
      W_myptr7_1405_delayed_8_0_1411_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr7_1405_delayed_8_0_1411_inst_req_1;
      W_myptr7_1405_delayed_8_0_1411_inst_ack_1<= rack(0);
      W_myptr7_1405_delayed_8_0_1411_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr7_1405_delayed_8_0_1411_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr7_1410,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr7_1405_delayed_8_0_1413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_myptr8_1428_delayed_8_0_1437_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_myptr8_1428_delayed_8_0_1437_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:W_myptr8_1428_delayed_8_0_1437_inst:started:   inputs: " & " myptr8_1436 = "& Convert_SLV_To_Hex_String(myptr8_1436));
          --
        end if; 
        if W_myptr8_1428_delayed_8_0_1437_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:W_myptr8_1428_delayed_8_0_1437_inst:finished:  outputs: " & " myptr8_1428_delayed_8_0_1439= "  & Convert_SLV_To_Hex_String(myptr8_1428_delayed_8_0_1439));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_myptr8_1428_delayed_8_0_1437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr8_1428_delayed_8_0_1437_inst_req_0;
      W_myptr8_1428_delayed_8_0_1437_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr8_1428_delayed_8_0_1437_inst_req_1;
      W_myptr8_1428_delayed_8_0_1437_inst_ack_1<= rack(0);
      W_myptr8_1428_delayed_8_0_1437_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr8_1428_delayed_8_0_1437_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr8_1436,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr8_1428_delayed_8_0_1439,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_1357_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_1357_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_1357_final_reg:started:   inputs: " & " array_obj_ref_1356_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1356_root_address));
          --
        end if; 
        if addr_of_1357_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_1357_final_reg:finished:  outputs: " & " myptr5_1358= "  & Convert_SLV_To_Hex_String(myptr5_1358));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_1357_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1357_final_reg_req_0;
      addr_of_1357_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1357_final_reg_req_1;
      addr_of_1357_final_reg_ack_1<= rack(0);
      addr_of_1357_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1357_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1356_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr5_1358,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_1383_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_1383_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_1383_final_reg:started:   inputs: " & " array_obj_ref_1382_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1382_root_address));
          --
        end if; 
        if addr_of_1383_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_1383_final_reg:finished:  outputs: " & " myptr6_1384= "  & Convert_SLV_To_Hex_String(myptr6_1384));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_1383_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1383_final_reg_req_0;
      addr_of_1383_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1383_final_reg_req_1;
      addr_of_1383_final_reg_ack_1<= rack(0);
      addr_of_1383_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1383_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1382_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr6_1384,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_1409_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_1409_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_1409_final_reg:started:   inputs: " & " array_obj_ref_1408_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1408_root_address));
          --
        end if; 
        if addr_of_1409_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_1409_final_reg:finished:  outputs: " & " myptr7_1410= "  & Convert_SLV_To_Hex_String(myptr7_1410));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_1409_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1409_final_reg_req_0;
      addr_of_1409_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1409_final_reg_req_1;
      addr_of_1409_final_reg_ack_1<= rack(0);
      addr_of_1409_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1409_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1408_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr7_1410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_1435_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_1435_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_1435_final_reg:started:   inputs: " & " array_obj_ref_1434_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1434_root_address));
          --
        end if; 
        if addr_of_1435_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_1435_final_reg:finished:  outputs: " & " myptr8_1436= "  & Convert_SLV_To_Hex_String(myptr8_1436));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_1435_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1435_final_reg_req_0;
      addr_of_1435_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1435_final_reg_req_1;
      addr_of_1435_final_reg_ack_1<= rack(0);
      addr_of_1435_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1435_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1434_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr8_1436,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_416_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_416_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_416_final_reg:started:   inputs: " & " array_obj_ref_415_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_415_root_address));
          --
        end if; 
        if addr_of_416_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_416_final_reg:finished:  outputs: " & " myptr1_417= "  & Convert_SLV_To_Hex_String(myptr1_417));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_416_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_416_final_reg_req_0;
      addr_of_416_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_416_final_reg_req_1;
      addr_of_416_final_reg_ack_1<= rack(0);
      addr_of_416_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_416_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_415_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr1_417,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_423_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_423_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_423_final_reg:started:   inputs: " & " array_obj_ref_422_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_422_root_address));
          --
        end if; 
        if addr_of_423_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_423_final_reg:finished:  outputs: " & " myptr2_424= "  & Convert_SLV_To_Hex_String(myptr2_424));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_423_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_423_final_reg_req_0;
      addr_of_423_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_423_final_reg_req_1;
      addr_of_423_final_reg_ack_1<= rack(0);
      addr_of_423_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_423_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_422_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr2_424,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_430_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_430_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_430_final_reg:started:   inputs: " & " array_obj_ref_429_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_429_root_address));
          --
        end if; 
        if addr_of_430_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_430_final_reg:finished:  outputs: " & " myptr3_431= "  & Convert_SLV_To_Hex_String(myptr3_431));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_430_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_430_final_reg_req_0;
      addr_of_430_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_430_final_reg_req_1;
      addr_of_430_final_reg_ack_1<= rack(0);
      addr_of_430_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_430_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_429_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr3_431,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_437_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_437_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_437_final_reg:started:   inputs: " & " array_obj_ref_436_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_436_root_address));
          --
        end if; 
        if addr_of_437_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:addr_of_437_final_reg:finished:  outputs: " & " myptr4_438= "  & Convert_SLV_To_Hex_String(myptr4_438));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_437_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_437_final_reg_req_0;
      addr_of_437_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_437_final_reg_req_1;
      addr_of_437_final_reg_ack_1<= rack(0);
      addr_of_437_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_437_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_436_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr4_438,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1365_inst flow-through 
    process(type_cast_1365_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1365_inst:flowthrough inputs: " & " out1_991 = "& Convert_SLV_To_Hex_String(out1_991) & " outputs:" & " type_cast_1365_wire= "  & Convert_SLV_To_Hex_String(type_cast_1365_wire));
      --
    end process; 
    -- interlock type_cast_1365_inst
    process(out1_991) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out1_991(15 downto 0);
      type_cast_1365_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1367_inst flow-through 
    process(type_cast_1367_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1367_inst:flowthrough inputs: " & " out2_1015 = "& Convert_SLV_To_Hex_String(out2_1015) & " outputs:" & " type_cast_1367_wire= "  & Convert_SLV_To_Hex_String(type_cast_1367_wire));
      --
    end process; 
    -- interlock type_cast_1367_inst
    process(out2_1015) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out2_1015(15 downto 0);
      type_cast_1367_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1370_inst flow-through 
    process(type_cast_1370_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1370_inst:flowthrough inputs: " & " out3_1039 = "& Convert_SLV_To_Hex_String(out3_1039) & " outputs:" & " type_cast_1370_wire= "  & Convert_SLV_To_Hex_String(type_cast_1370_wire));
      --
    end process; 
    -- interlock type_cast_1370_inst
    process(out3_1039) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out3_1039(15 downto 0);
      type_cast_1370_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1372_inst flow-through 
    process(type_cast_1372_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1372_inst:flowthrough inputs: " & " out4_1063 = "& Convert_SLV_To_Hex_String(out4_1063) & " outputs:" & " type_cast_1372_wire= "  & Convert_SLV_To_Hex_String(type_cast_1372_wire));
      --
    end process; 
    -- interlock type_cast_1372_inst
    process(out4_1063) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out4_1063(15 downto 0);
      type_cast_1372_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1391_inst flow-through 
    process(type_cast_1391_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1391_inst:flowthrough inputs: " & " out5_1087 = "& Convert_SLV_To_Hex_String(out5_1087) & " outputs:" & " type_cast_1391_wire= "  & Convert_SLV_To_Hex_String(type_cast_1391_wire));
      --
    end process; 
    -- interlock type_cast_1391_inst
    process(out5_1087) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out5_1087(15 downto 0);
      type_cast_1391_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1393_inst flow-through 
    process(type_cast_1393_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1393_inst:flowthrough inputs: " & " out6_1111 = "& Convert_SLV_To_Hex_String(out6_1111) & " outputs:" & " type_cast_1393_wire= "  & Convert_SLV_To_Hex_String(type_cast_1393_wire));
      --
    end process; 
    -- interlock type_cast_1393_inst
    process(out6_1111) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out6_1111(15 downto 0);
      type_cast_1393_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1396_inst flow-through 
    process(type_cast_1396_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1396_inst:flowthrough inputs: " & " out7_1135 = "& Convert_SLV_To_Hex_String(out7_1135) & " outputs:" & " type_cast_1396_wire= "  & Convert_SLV_To_Hex_String(type_cast_1396_wire));
      --
    end process; 
    -- interlock type_cast_1396_inst
    process(out7_1135) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out7_1135(15 downto 0);
      type_cast_1396_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1398_inst flow-through 
    process(type_cast_1398_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1398_inst:flowthrough inputs: " & " out8_1159 = "& Convert_SLV_To_Hex_String(out8_1159) & " outputs:" & " type_cast_1398_wire= "  & Convert_SLV_To_Hex_String(type_cast_1398_wire));
      --
    end process; 
    -- interlock type_cast_1398_inst
    process(out8_1159) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out8_1159(15 downto 0);
      type_cast_1398_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1417_inst flow-through 
    process(type_cast_1417_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1417_inst:flowthrough inputs: " & " out9_1183 = "& Convert_SLV_To_Hex_String(out9_1183) & " outputs:" & " type_cast_1417_wire= "  & Convert_SLV_To_Hex_String(type_cast_1417_wire));
      --
    end process; 
    -- interlock type_cast_1417_inst
    process(out9_1183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out9_1183(15 downto 0);
      type_cast_1417_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1419_inst flow-through 
    process(type_cast_1419_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1419_inst:flowthrough inputs: " & " out10_1207 = "& Convert_SLV_To_Hex_String(out10_1207) & " outputs:" & " type_cast_1419_wire= "  & Convert_SLV_To_Hex_String(type_cast_1419_wire));
      --
    end process; 
    -- interlock type_cast_1419_inst
    process(out10_1207) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out10_1207(15 downto 0);
      type_cast_1419_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1422_inst flow-through 
    process(type_cast_1422_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1422_inst:flowthrough inputs: " & " out11_1231 = "& Convert_SLV_To_Hex_String(out11_1231) & " outputs:" & " type_cast_1422_wire= "  & Convert_SLV_To_Hex_String(type_cast_1422_wire));
      --
    end process; 
    -- interlock type_cast_1422_inst
    process(out11_1231) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out11_1231(15 downto 0);
      type_cast_1422_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1424_inst flow-through 
    process(type_cast_1424_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1424_inst:flowthrough inputs: " & " out12_1255 = "& Convert_SLV_To_Hex_String(out12_1255) & " outputs:" & " type_cast_1424_wire= "  & Convert_SLV_To_Hex_String(type_cast_1424_wire));
      --
    end process; 
    -- interlock type_cast_1424_inst
    process(out12_1255) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out12_1255(15 downto 0);
      type_cast_1424_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1443_inst flow-through 
    process(type_cast_1443_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1443_inst:flowthrough inputs: " & " out13_1279 = "& Convert_SLV_To_Hex_String(out13_1279) & " outputs:" & " type_cast_1443_wire= "  & Convert_SLV_To_Hex_String(type_cast_1443_wire));
      --
    end process; 
    -- interlock type_cast_1443_inst
    process(out13_1279) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out13_1279(15 downto 0);
      type_cast_1443_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1445_inst flow-through 
    process(type_cast_1445_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1445_inst:flowthrough inputs: " & " out14_1303 = "& Convert_SLV_To_Hex_String(out14_1303) & " outputs:" & " type_cast_1445_wire= "  & Convert_SLV_To_Hex_String(type_cast_1445_wire));
      --
    end process; 
    -- interlock type_cast_1445_inst
    process(out14_1303) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out14_1303(15 downto 0);
      type_cast_1445_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1448_inst flow-through 
    process(type_cast_1448_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1448_inst:flowthrough inputs: " & " out15_1327 = "& Convert_SLV_To_Hex_String(out15_1327) & " outputs:" & " type_cast_1448_wire= "  & Convert_SLV_To_Hex_String(type_cast_1448_wire));
      --
    end process; 
    -- interlock type_cast_1448_inst
    process(out15_1327) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out15_1327(15 downto 0);
      type_cast_1448_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1450_inst flow-through 
    process(type_cast_1450_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1450_inst:flowthrough inputs: " & " out16_1351 = "& Convert_SLV_To_Hex_String(out16_1351) & " outputs:" & " type_cast_1450_wire= "  & Convert_SLV_To_Hex_String(type_cast_1450_wire));
      --
    end process; 
    -- interlock type_cast_1450_inst
    process(out16_1351) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out16_1351(15 downto 0);
      type_cast_1450_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1456_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1456_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1456_inst:started:   inputs: " & " out1_991 = "& Convert_SLV_To_Hex_String(out1_991));
          --
        end if; 
        if type_cast_1456_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_1456_inst:finished:  outputs: " & " output_buffer= "  & Convert_SLV_To_Hex_String(output_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1456_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1456_inst_req_0;
      type_cast_1456_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1456_inst_req_1;
      type_cast_1456_inst_ack_1<= rack(0);
      type_cast_1456_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1456_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => out1_991,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_714_inst flow-through 
    process(a11_715) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_714_inst:flowthrough inputs: " & " sliced_v11_458 = "& Convert_SLV_To_Hex_String(sliced_v11_458) & " outputs:" & " a11_715= "  & Convert_SLV_To_Hex_String(a11_715));
      --
    end process; 
    -- interlock type_cast_714_inst
    process(sliced_v11_458) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v11_458(15 downto 0);
      a11_715 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_718_inst flow-through 
    process(a12_719) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_718_inst:flowthrough inputs: " & " sliced_v12_462 = "& Convert_SLV_To_Hex_String(sliced_v12_462) & " outputs:" & " a12_719= "  & Convert_SLV_To_Hex_String(a12_719));
      --
    end process; 
    -- interlock type_cast_718_inst
    process(sliced_v12_462) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v12_462(15 downto 0);
      a12_719 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_722_inst flow-through 
    process(a13_723) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_722_inst:flowthrough inputs: " & " sliced_v13_466 = "& Convert_SLV_To_Hex_String(sliced_v13_466) & " outputs:" & " a13_723= "  & Convert_SLV_To_Hex_String(a13_723));
      --
    end process; 
    -- interlock type_cast_722_inst
    process(sliced_v13_466) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v13_466(15 downto 0);
      a13_723 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_726_inst flow-through 
    process(a14_727) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_726_inst:flowthrough inputs: " & " sliced_v14_470 = "& Convert_SLV_To_Hex_String(sliced_v14_470) & " outputs:" & " a14_727= "  & Convert_SLV_To_Hex_String(a14_727));
      --
    end process; 
    -- interlock type_cast_726_inst
    process(sliced_v14_470) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v14_470(15 downto 0);
      a14_727 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_730_inst flow-through 
    process(a15_731) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_730_inst:flowthrough inputs: " & " sliced_v15_474 = "& Convert_SLV_To_Hex_String(sliced_v15_474) & " outputs:" & " a15_731= "  & Convert_SLV_To_Hex_String(a15_731));
      --
    end process; 
    -- interlock type_cast_730_inst
    process(sliced_v15_474) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v15_474(15 downto 0);
      a15_731 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_734_inst flow-through 
    process(a16_735) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_734_inst:flowthrough inputs: " & " sliced_v16_478 = "& Convert_SLV_To_Hex_String(sliced_v16_478) & " outputs:" & " a16_735= "  & Convert_SLV_To_Hex_String(a16_735));
      --
    end process; 
    -- interlock type_cast_734_inst
    process(sliced_v16_478) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v16_478(15 downto 0);
      a16_735 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_738_inst flow-through 
    process(a17_739) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_738_inst:flowthrough inputs: " & " sliced_v17_482 = "& Convert_SLV_To_Hex_String(sliced_v17_482) & " outputs:" & " a17_739= "  & Convert_SLV_To_Hex_String(a17_739));
      --
    end process; 
    -- interlock type_cast_738_inst
    process(sliced_v17_482) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v17_482(15 downto 0);
      a17_739 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_742_inst flow-through 
    process(a18_743) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_742_inst:flowthrough inputs: " & " sliced_v18_486 = "& Convert_SLV_To_Hex_String(sliced_v18_486) & " outputs:" & " a18_743= "  & Convert_SLV_To_Hex_String(a18_743));
      --
    end process; 
    -- interlock type_cast_742_inst
    process(sliced_v18_486) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v18_486(15 downto 0);
      a18_743 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_746_inst flow-through 
    process(a19_747) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_746_inst:flowthrough inputs: " & " sliced_v19_490 = "& Convert_SLV_To_Hex_String(sliced_v19_490) & " outputs:" & " a19_747= "  & Convert_SLV_To_Hex_String(a19_747));
      --
    end process; 
    -- interlock type_cast_746_inst
    process(sliced_v19_490) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v19_490(15 downto 0);
      a19_747 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_750_inst flow-through 
    process(a110_751) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_750_inst:flowthrough inputs: " & " sliced_v110_494 = "& Convert_SLV_To_Hex_String(sliced_v110_494) & " outputs:" & " a110_751= "  & Convert_SLV_To_Hex_String(a110_751));
      --
    end process; 
    -- interlock type_cast_750_inst
    process(sliced_v110_494) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v110_494(15 downto 0);
      a110_751 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_754_inst flow-through 
    process(a111_755) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_754_inst:flowthrough inputs: " & " sliced_v111_498 = "& Convert_SLV_To_Hex_String(sliced_v111_498) & " outputs:" & " a111_755= "  & Convert_SLV_To_Hex_String(a111_755));
      --
    end process; 
    -- interlock type_cast_754_inst
    process(sliced_v111_498) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v111_498(15 downto 0);
      a111_755 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_758_inst flow-through 
    process(a112_759) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_758_inst:flowthrough inputs: " & " sliced_v112_502 = "& Convert_SLV_To_Hex_String(sliced_v112_502) & " outputs:" & " a112_759= "  & Convert_SLV_To_Hex_String(a112_759));
      --
    end process; 
    -- interlock type_cast_758_inst
    process(sliced_v112_502) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v112_502(15 downto 0);
      a112_759 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_762_inst flow-through 
    process(a113_763) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_762_inst:flowthrough inputs: " & " sliced_v113_506 = "& Convert_SLV_To_Hex_String(sliced_v113_506) & " outputs:" & " a113_763= "  & Convert_SLV_To_Hex_String(a113_763));
      --
    end process; 
    -- interlock type_cast_762_inst
    process(sliced_v113_506) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v113_506(15 downto 0);
      a113_763 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_766_inst flow-through 
    process(a114_767) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_766_inst:flowthrough inputs: " & " sliced_v114_510 = "& Convert_SLV_To_Hex_String(sliced_v114_510) & " outputs:" & " a114_767= "  & Convert_SLV_To_Hex_String(a114_767));
      --
    end process; 
    -- interlock type_cast_766_inst
    process(sliced_v114_510) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v114_510(15 downto 0);
      a114_767 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_770_inst flow-through 
    process(a115_771) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_770_inst:flowthrough inputs: " & " sliced_v115_514 = "& Convert_SLV_To_Hex_String(sliced_v115_514) & " outputs:" & " a115_771= "  & Convert_SLV_To_Hex_String(a115_771));
      --
    end process; 
    -- interlock type_cast_770_inst
    process(sliced_v115_514) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v115_514(15 downto 0);
      a115_771 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_774_inst flow-through 
    process(a116_775) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_774_inst:flowthrough inputs: " & " sliced_v116_518 = "& Convert_SLV_To_Hex_String(sliced_v116_518) & " outputs:" & " a116_775= "  & Convert_SLV_To_Hex_String(a116_775));
      --
    end process; 
    -- interlock type_cast_774_inst
    process(sliced_v116_518) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v116_518(15 downto 0);
      a116_775 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_778_inst flow-through 
    process(a21_779) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_778_inst:flowthrough inputs: " & " sliced_v21_522 = "& Convert_SLV_To_Hex_String(sliced_v21_522) & " outputs:" & " a21_779= "  & Convert_SLV_To_Hex_String(a21_779));
      --
    end process; 
    -- interlock type_cast_778_inst
    process(sliced_v21_522) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v21_522(15 downto 0);
      a21_779 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_782_inst flow-through 
    process(a22_783) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_782_inst:flowthrough inputs: " & " sliced_v22_526 = "& Convert_SLV_To_Hex_String(sliced_v22_526) & " outputs:" & " a22_783= "  & Convert_SLV_To_Hex_String(a22_783));
      --
    end process; 
    -- interlock type_cast_782_inst
    process(sliced_v22_526) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v22_526(15 downto 0);
      a22_783 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_786_inst flow-through 
    process(a23_787) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_786_inst:flowthrough inputs: " & " sliced_v23_530 = "& Convert_SLV_To_Hex_String(sliced_v23_530) & " outputs:" & " a23_787= "  & Convert_SLV_To_Hex_String(a23_787));
      --
    end process; 
    -- interlock type_cast_786_inst
    process(sliced_v23_530) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v23_530(15 downto 0);
      a23_787 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_790_inst flow-through 
    process(a24_791) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_790_inst:flowthrough inputs: " & " sliced_v24_534 = "& Convert_SLV_To_Hex_String(sliced_v24_534) & " outputs:" & " a24_791= "  & Convert_SLV_To_Hex_String(a24_791));
      --
    end process; 
    -- interlock type_cast_790_inst
    process(sliced_v24_534) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v24_534(15 downto 0);
      a24_791 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_794_inst flow-through 
    process(a25_795) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_794_inst:flowthrough inputs: " & " sliced_v25_538 = "& Convert_SLV_To_Hex_String(sliced_v25_538) & " outputs:" & " a25_795= "  & Convert_SLV_To_Hex_String(a25_795));
      --
    end process; 
    -- interlock type_cast_794_inst
    process(sliced_v25_538) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v25_538(15 downto 0);
      a25_795 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_798_inst flow-through 
    process(a26_799) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_798_inst:flowthrough inputs: " & " sliced_v26_542 = "& Convert_SLV_To_Hex_String(sliced_v26_542) & " outputs:" & " a26_799= "  & Convert_SLV_To_Hex_String(a26_799));
      --
    end process; 
    -- interlock type_cast_798_inst
    process(sliced_v26_542) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v26_542(15 downto 0);
      a26_799 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_802_inst flow-through 
    process(a27_803) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_802_inst:flowthrough inputs: " & " sliced_v27_546 = "& Convert_SLV_To_Hex_String(sliced_v27_546) & " outputs:" & " a27_803= "  & Convert_SLV_To_Hex_String(a27_803));
      --
    end process; 
    -- interlock type_cast_802_inst
    process(sliced_v27_546) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v27_546(15 downto 0);
      a27_803 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_806_inst flow-through 
    process(a28_807) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_806_inst:flowthrough inputs: " & " sliced_v28_550 = "& Convert_SLV_To_Hex_String(sliced_v28_550) & " outputs:" & " a28_807= "  & Convert_SLV_To_Hex_String(a28_807));
      --
    end process; 
    -- interlock type_cast_806_inst
    process(sliced_v28_550) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v28_550(15 downto 0);
      a28_807 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_810_inst flow-through 
    process(a29_811) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_810_inst:flowthrough inputs: " & " sliced_v29_554 = "& Convert_SLV_To_Hex_String(sliced_v29_554) & " outputs:" & " a29_811= "  & Convert_SLV_To_Hex_String(a29_811));
      --
    end process; 
    -- interlock type_cast_810_inst
    process(sliced_v29_554) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v29_554(15 downto 0);
      a29_811 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_814_inst flow-through 
    process(a210_815) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_814_inst:flowthrough inputs: " & " sliced_v210_558 = "& Convert_SLV_To_Hex_String(sliced_v210_558) & " outputs:" & " a210_815= "  & Convert_SLV_To_Hex_String(a210_815));
      --
    end process; 
    -- interlock type_cast_814_inst
    process(sliced_v210_558) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v210_558(15 downto 0);
      a210_815 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_818_inst flow-through 
    process(a211_819) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_818_inst:flowthrough inputs: " & " sliced_v211_562 = "& Convert_SLV_To_Hex_String(sliced_v211_562) & " outputs:" & " a211_819= "  & Convert_SLV_To_Hex_String(a211_819));
      --
    end process; 
    -- interlock type_cast_818_inst
    process(sliced_v211_562) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v211_562(15 downto 0);
      a211_819 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_822_inst flow-through 
    process(a212_823) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_822_inst:flowthrough inputs: " & " sliced_v212_566 = "& Convert_SLV_To_Hex_String(sliced_v212_566) & " outputs:" & " a212_823= "  & Convert_SLV_To_Hex_String(a212_823));
      --
    end process; 
    -- interlock type_cast_822_inst
    process(sliced_v212_566) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v212_566(15 downto 0);
      a212_823 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_826_inst flow-through 
    process(a213_827) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_826_inst:flowthrough inputs: " & " sliced_v213_570 = "& Convert_SLV_To_Hex_String(sliced_v213_570) & " outputs:" & " a213_827= "  & Convert_SLV_To_Hex_String(a213_827));
      --
    end process; 
    -- interlock type_cast_826_inst
    process(sliced_v213_570) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v213_570(15 downto 0);
      a213_827 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_830_inst flow-through 
    process(a214_831) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_830_inst:flowthrough inputs: " & " sliced_v214_574 = "& Convert_SLV_To_Hex_String(sliced_v214_574) & " outputs:" & " a214_831= "  & Convert_SLV_To_Hex_String(a214_831));
      --
    end process; 
    -- interlock type_cast_830_inst
    process(sliced_v214_574) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v214_574(15 downto 0);
      a214_831 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_834_inst flow-through 
    process(a215_835) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_834_inst:flowthrough inputs: " & " sliced_v215_578 = "& Convert_SLV_To_Hex_String(sliced_v215_578) & " outputs:" & " a215_835= "  & Convert_SLV_To_Hex_String(a215_835));
      --
    end process; 
    -- interlock type_cast_834_inst
    process(sliced_v215_578) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v215_578(15 downto 0);
      a215_835 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_838_inst flow-through 
    process(a216_839) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_838_inst:flowthrough inputs: " & " sliced_v216_582 = "& Convert_SLV_To_Hex_String(sliced_v216_582) & " outputs:" & " a216_839= "  & Convert_SLV_To_Hex_String(a216_839));
      --
    end process; 
    -- interlock type_cast_838_inst
    process(sliced_v216_582) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v216_582(15 downto 0);
      a216_839 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_842_inst flow-through 
    process(a31_843) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_842_inst:flowthrough inputs: " & " sliced_v31_586 = "& Convert_SLV_To_Hex_String(sliced_v31_586) & " outputs:" & " a31_843= "  & Convert_SLV_To_Hex_String(a31_843));
      --
    end process; 
    -- interlock type_cast_842_inst
    process(sliced_v31_586) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v31_586(15 downto 0);
      a31_843 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_846_inst flow-through 
    process(a32_847) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_846_inst:flowthrough inputs: " & " sliced_v32_590 = "& Convert_SLV_To_Hex_String(sliced_v32_590) & " outputs:" & " a32_847= "  & Convert_SLV_To_Hex_String(a32_847));
      --
    end process; 
    -- interlock type_cast_846_inst
    process(sliced_v32_590) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v32_590(15 downto 0);
      a32_847 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_850_inst flow-through 
    process(a33_851) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_850_inst:flowthrough inputs: " & " sliced_v33_594 = "& Convert_SLV_To_Hex_String(sliced_v33_594) & " outputs:" & " a33_851= "  & Convert_SLV_To_Hex_String(a33_851));
      --
    end process; 
    -- interlock type_cast_850_inst
    process(sliced_v33_594) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v33_594(15 downto 0);
      a33_851 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_854_inst flow-through 
    process(a34_855) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_854_inst:flowthrough inputs: " & " sliced_v34_598 = "& Convert_SLV_To_Hex_String(sliced_v34_598) & " outputs:" & " a34_855= "  & Convert_SLV_To_Hex_String(a34_855));
      --
    end process; 
    -- interlock type_cast_854_inst
    process(sliced_v34_598) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v34_598(15 downto 0);
      a34_855 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_858_inst flow-through 
    process(a35_859) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_858_inst:flowthrough inputs: " & " sliced_v35_602 = "& Convert_SLV_To_Hex_String(sliced_v35_602) & " outputs:" & " a35_859= "  & Convert_SLV_To_Hex_String(a35_859));
      --
    end process; 
    -- interlock type_cast_858_inst
    process(sliced_v35_602) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v35_602(15 downto 0);
      a35_859 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_862_inst flow-through 
    process(a36_863) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_862_inst:flowthrough inputs: " & " sliced_v36_606 = "& Convert_SLV_To_Hex_String(sliced_v36_606) & " outputs:" & " a36_863= "  & Convert_SLV_To_Hex_String(a36_863));
      --
    end process; 
    -- interlock type_cast_862_inst
    process(sliced_v36_606) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v36_606(15 downto 0);
      a36_863 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_866_inst flow-through 
    process(a37_867) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_866_inst:flowthrough inputs: " & " sliced_v37_610 = "& Convert_SLV_To_Hex_String(sliced_v37_610) & " outputs:" & " a37_867= "  & Convert_SLV_To_Hex_String(a37_867));
      --
    end process; 
    -- interlock type_cast_866_inst
    process(sliced_v37_610) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v37_610(15 downto 0);
      a37_867 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_870_inst flow-through 
    process(a38_871) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_870_inst:flowthrough inputs: " & " sliced_v38_614 = "& Convert_SLV_To_Hex_String(sliced_v38_614) & " outputs:" & " a38_871= "  & Convert_SLV_To_Hex_String(a38_871));
      --
    end process; 
    -- interlock type_cast_870_inst
    process(sliced_v38_614) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v38_614(15 downto 0);
      a38_871 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_874_inst flow-through 
    process(a39_875) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_874_inst:flowthrough inputs: " & " sliced_v39_618 = "& Convert_SLV_To_Hex_String(sliced_v39_618) & " outputs:" & " a39_875= "  & Convert_SLV_To_Hex_String(a39_875));
      --
    end process; 
    -- interlock type_cast_874_inst
    process(sliced_v39_618) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v39_618(15 downto 0);
      a39_875 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_878_inst flow-through 
    process(a310_879) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_878_inst:flowthrough inputs: " & " sliced_v310_622 = "& Convert_SLV_To_Hex_String(sliced_v310_622) & " outputs:" & " a310_879= "  & Convert_SLV_To_Hex_String(a310_879));
      --
    end process; 
    -- interlock type_cast_878_inst
    process(sliced_v310_622) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v310_622(15 downto 0);
      a310_879 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_882_inst flow-through 
    process(a311_883) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_882_inst:flowthrough inputs: " & " sliced_v311_626 = "& Convert_SLV_To_Hex_String(sliced_v311_626) & " outputs:" & " a311_883= "  & Convert_SLV_To_Hex_String(a311_883));
      --
    end process; 
    -- interlock type_cast_882_inst
    process(sliced_v311_626) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v311_626(15 downto 0);
      a311_883 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_886_inst flow-through 
    process(a312_887) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_886_inst:flowthrough inputs: " & " sliced_v312_630 = "& Convert_SLV_To_Hex_String(sliced_v312_630) & " outputs:" & " a312_887= "  & Convert_SLV_To_Hex_String(a312_887));
      --
    end process; 
    -- interlock type_cast_886_inst
    process(sliced_v312_630) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v312_630(15 downto 0);
      a312_887 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_890_inst flow-through 
    process(a313_891) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_890_inst:flowthrough inputs: " & " sliced_v313_634 = "& Convert_SLV_To_Hex_String(sliced_v313_634) & " outputs:" & " a313_891= "  & Convert_SLV_To_Hex_String(a313_891));
      --
    end process; 
    -- interlock type_cast_890_inst
    process(sliced_v313_634) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v313_634(15 downto 0);
      a313_891 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_894_inst flow-through 
    process(a314_895) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_894_inst:flowthrough inputs: " & " sliced_v314_638 = "& Convert_SLV_To_Hex_String(sliced_v314_638) & " outputs:" & " a314_895= "  & Convert_SLV_To_Hex_String(a314_895));
      --
    end process; 
    -- interlock type_cast_894_inst
    process(sliced_v314_638) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v314_638(15 downto 0);
      a314_895 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_898_inst flow-through 
    process(a315_899) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_898_inst:flowthrough inputs: " & " sliced_v315_642 = "& Convert_SLV_To_Hex_String(sliced_v315_642) & " outputs:" & " a315_899= "  & Convert_SLV_To_Hex_String(a315_899));
      --
    end process; 
    -- interlock type_cast_898_inst
    process(sliced_v315_642) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v315_642(15 downto 0);
      a315_899 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_902_inst flow-through 
    process(a316_903) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_902_inst:flowthrough inputs: " & " sliced_v316_646 = "& Convert_SLV_To_Hex_String(sliced_v316_646) & " outputs:" & " a316_903= "  & Convert_SLV_To_Hex_String(a316_903));
      --
    end process; 
    -- interlock type_cast_902_inst
    process(sliced_v316_646) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v316_646(15 downto 0);
      a316_903 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_906_inst flow-through 
    process(a41_907) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_906_inst:flowthrough inputs: " & " sliced_v41_650 = "& Convert_SLV_To_Hex_String(sliced_v41_650) & " outputs:" & " a41_907= "  & Convert_SLV_To_Hex_String(a41_907));
      --
    end process; 
    -- interlock type_cast_906_inst
    process(sliced_v41_650) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v41_650(15 downto 0);
      a41_907 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_910_inst flow-through 
    process(a42_911) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_910_inst:flowthrough inputs: " & " sliced_v42_654 = "& Convert_SLV_To_Hex_String(sliced_v42_654) & " outputs:" & " a42_911= "  & Convert_SLV_To_Hex_String(a42_911));
      --
    end process; 
    -- interlock type_cast_910_inst
    process(sliced_v42_654) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v42_654(15 downto 0);
      a42_911 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_914_inst flow-through 
    process(a43_915) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_914_inst:flowthrough inputs: " & " sliced_v43_658 = "& Convert_SLV_To_Hex_String(sliced_v43_658) & " outputs:" & " a43_915= "  & Convert_SLV_To_Hex_String(a43_915));
      --
    end process; 
    -- interlock type_cast_914_inst
    process(sliced_v43_658) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v43_658(15 downto 0);
      a43_915 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_918_inst flow-through 
    process(a44_919) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_918_inst:flowthrough inputs: " & " sliced_v44_662 = "& Convert_SLV_To_Hex_String(sliced_v44_662) & " outputs:" & " a44_919= "  & Convert_SLV_To_Hex_String(a44_919));
      --
    end process; 
    -- interlock type_cast_918_inst
    process(sliced_v44_662) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v44_662(15 downto 0);
      a44_919 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_922_inst flow-through 
    process(a45_923) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_922_inst:flowthrough inputs: " & " sliced_v45_666 = "& Convert_SLV_To_Hex_String(sliced_v45_666) & " outputs:" & " a45_923= "  & Convert_SLV_To_Hex_String(a45_923));
      --
    end process; 
    -- interlock type_cast_922_inst
    process(sliced_v45_666) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v45_666(15 downto 0);
      a45_923 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_926_inst flow-through 
    process(a46_927) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_926_inst:flowthrough inputs: " & " sliced_v46_670 = "& Convert_SLV_To_Hex_String(sliced_v46_670) & " outputs:" & " a46_927= "  & Convert_SLV_To_Hex_String(a46_927));
      --
    end process; 
    -- interlock type_cast_926_inst
    process(sliced_v46_670) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v46_670(15 downto 0);
      a46_927 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_930_inst flow-through 
    process(a47_931) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_930_inst:flowthrough inputs: " & " sliced_v47_674 = "& Convert_SLV_To_Hex_String(sliced_v47_674) & " outputs:" & " a47_931= "  & Convert_SLV_To_Hex_String(a47_931));
      --
    end process; 
    -- interlock type_cast_930_inst
    process(sliced_v47_674) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v47_674(15 downto 0);
      a47_931 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_934_inst flow-through 
    process(a48_935) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_934_inst:flowthrough inputs: " & " sliced_v48_678 = "& Convert_SLV_To_Hex_String(sliced_v48_678) & " outputs:" & " a48_935= "  & Convert_SLV_To_Hex_String(a48_935));
      --
    end process; 
    -- interlock type_cast_934_inst
    process(sliced_v48_678) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v48_678(15 downto 0);
      a48_935 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_938_inst flow-through 
    process(a49_939) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_938_inst:flowthrough inputs: " & " sliced_v49_682 = "& Convert_SLV_To_Hex_String(sliced_v49_682) & " outputs:" & " a49_939= "  & Convert_SLV_To_Hex_String(a49_939));
      --
    end process; 
    -- interlock type_cast_938_inst
    process(sliced_v49_682) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v49_682(15 downto 0);
      a49_939 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_942_inst flow-through 
    process(a410_943) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_942_inst:flowthrough inputs: " & " sliced_v410_686 = "& Convert_SLV_To_Hex_String(sliced_v410_686) & " outputs:" & " a410_943= "  & Convert_SLV_To_Hex_String(a410_943));
      --
    end process; 
    -- interlock type_cast_942_inst
    process(sliced_v410_686) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v410_686(15 downto 0);
      a410_943 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_946_inst flow-through 
    process(a411_947) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_946_inst:flowthrough inputs: " & " sliced_v411_690 = "& Convert_SLV_To_Hex_String(sliced_v411_690) & " outputs:" & " a411_947= "  & Convert_SLV_To_Hex_String(a411_947));
      --
    end process; 
    -- interlock type_cast_946_inst
    process(sliced_v411_690) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v411_690(15 downto 0);
      a411_947 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_950_inst flow-through 
    process(a412_951) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_950_inst:flowthrough inputs: " & " sliced_v412_694 = "& Convert_SLV_To_Hex_String(sliced_v412_694) & " outputs:" & " a412_951= "  & Convert_SLV_To_Hex_String(a412_951));
      --
    end process; 
    -- interlock type_cast_950_inst
    process(sliced_v412_694) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v412_694(15 downto 0);
      a412_951 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_954_inst flow-through 
    process(a413_955) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_954_inst:flowthrough inputs: " & " sliced_v413_698 = "& Convert_SLV_To_Hex_String(sliced_v413_698) & " outputs:" & " a413_955= "  & Convert_SLV_To_Hex_String(a413_955));
      --
    end process; 
    -- interlock type_cast_954_inst
    process(sliced_v413_698) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v413_698(15 downto 0);
      a413_955 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_958_inst flow-through 
    process(a414_959) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_958_inst:flowthrough inputs: " & " sliced_v414_702 = "& Convert_SLV_To_Hex_String(sliced_v414_702) & " outputs:" & " a414_959= "  & Convert_SLV_To_Hex_String(a414_959));
      --
    end process; 
    -- interlock type_cast_958_inst
    process(sliced_v414_702) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v414_702(15 downto 0);
      a414_959 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_962_inst flow-through 
    process(a415_963) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_962_inst:flowthrough inputs: " & " sliced_v415_706 = "& Convert_SLV_To_Hex_String(sliced_v415_706) & " outputs:" & " a415_963= "  & Convert_SLV_To_Hex_String(a415_963));
      --
    end process; 
    -- interlock type_cast_962_inst
    process(sliced_v415_706) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v415_706(15 downto 0);
      a415_963 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_966_inst flow-through 
    process(a416_967) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:type_cast_966_inst:flowthrough inputs: " & " sliced_v416_710 = "& Convert_SLV_To_Hex_String(sliced_v416_710) & " outputs:" & " a416_967= "  & Convert_SLV_To_Hex_String(a416_967));
      --
    end process; 
    -- interlock type_cast_966_inst
    process(sliced_v416_710) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v416_710(15 downto 0);
      a416_967 <= tmp_var; -- 
    end process;
    -- logger for operator array_obj_ref_1356_index_1_rename flow-through 
    process(R_addr_1355_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1356_index_1_rename:flowthrough  inputs: " & " R_addr_1355_resized = "& Convert_SLV_To_Hex_String(R_addr_1355_resized) & "outputs: " & " R_addr_1355_scaled= "  & Convert_SLV_To_Hex_String(R_addr_1355_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1356_index_1_rename
    process(R_addr_1355_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_1355_resized;
      ov(13 downto 0) := iv;
      R_addr_1355_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1356_index_1_resize flow-through 
    process(R_addr_1355_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1356_index_1_resize:flowthrough  inputs: " & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & "outputs: " & " R_addr_1355_resized= "  & Convert_SLV_To_Hex_String(R_addr_1355_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1356_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(13 downto 0);
      R_addr_1355_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1356_root_address_inst flow-through 
    process(array_obj_ref_1356_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1356_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1356_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1356_final_offset) & "outputs: " & " array_obj_ref_1356_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1356_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1356_root_address_inst
    process(array_obj_ref_1356_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1356_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1356_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1382_index_1_rename flow-through 
    process(ADD_u32_u32_1381_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1382_index_1_rename:flowthrough  inputs: " & " ADD_u32_u32_1381_resized = "& Convert_SLV_To_Hex_String(ADD_u32_u32_1381_resized) & "outputs: " & " ADD_u32_u32_1381_scaled= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_1381_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1382_index_1_rename
    process(ADD_u32_u32_1381_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1381_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1381_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1382_index_1_resize flow-through 
    process(ADD_u32_u32_1381_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1382_index_1_resize:flowthrough  inputs: " & " ADD_u32_u32_1381_wire = "& Convert_SLV_To_Hex_String(ADD_u32_u32_1381_wire) & "outputs: " & " ADD_u32_u32_1381_resized= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_1381_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1382_index_1_resize
    process(ADD_u32_u32_1381_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1381_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1381_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1382_root_address_inst flow-through 
    process(array_obj_ref_1382_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1382_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1382_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1382_final_offset) & "outputs: " & " array_obj_ref_1382_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1382_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1382_root_address_inst
    process(array_obj_ref_1382_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1382_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1382_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1408_index_1_rename flow-through 
    process(ADD_u32_u32_1407_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1408_index_1_rename:flowthrough  inputs: " & " ADD_u32_u32_1407_resized = "& Convert_SLV_To_Hex_String(ADD_u32_u32_1407_resized) & "outputs: " & " ADD_u32_u32_1407_scaled= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_1407_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1408_index_1_rename
    process(ADD_u32_u32_1407_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1407_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1407_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1408_index_1_resize flow-through 
    process(ADD_u32_u32_1407_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1408_index_1_resize:flowthrough  inputs: " & " ADD_u32_u32_1407_wire = "& Convert_SLV_To_Hex_String(ADD_u32_u32_1407_wire) & "outputs: " & " ADD_u32_u32_1407_resized= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_1407_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1408_index_1_resize
    process(ADD_u32_u32_1407_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1407_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1407_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1408_root_address_inst flow-through 
    process(array_obj_ref_1408_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1408_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1408_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1408_final_offset) & "outputs: " & " array_obj_ref_1408_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1408_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1408_root_address_inst
    process(array_obj_ref_1408_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1408_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1408_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1434_index_1_rename flow-through 
    process(ADD_u32_u32_1433_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1434_index_1_rename:flowthrough  inputs: " & " ADD_u32_u32_1433_resized = "& Convert_SLV_To_Hex_String(ADD_u32_u32_1433_resized) & "outputs: " & " ADD_u32_u32_1433_scaled= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_1433_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1434_index_1_rename
    process(ADD_u32_u32_1433_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1433_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1433_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1434_index_1_resize flow-through 
    process(ADD_u32_u32_1433_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1434_index_1_resize:flowthrough  inputs: " & " ADD_u32_u32_1433_wire = "& Convert_SLV_To_Hex_String(ADD_u32_u32_1433_wire) & "outputs: " & " ADD_u32_u32_1433_resized= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_1433_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1434_index_1_resize
    process(ADD_u32_u32_1433_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1433_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1433_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1434_root_address_inst flow-through 
    process(array_obj_ref_1434_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1434_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1434_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1434_final_offset) & "outputs: " & " array_obj_ref_1434_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1434_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1434_root_address_inst
    process(array_obj_ref_1434_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1434_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1434_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_415_index_1_rename flow-through 
    process(R_addr1_414_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_415_index_1_rename:flowthrough  inputs: " & " R_addr1_414_resized = "& Convert_SLV_To_Hex_String(R_addr1_414_resized) & "outputs: " & " R_addr1_414_scaled= "  & Convert_SLV_To_Hex_String(R_addr1_414_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_415_index_1_rename
    process(R_addr1_414_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr1_414_resized;
      ov(13 downto 0) := iv;
      R_addr1_414_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_415_index_1_resize flow-through 
    process(R_addr1_414_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_415_index_1_resize:flowthrough  inputs: " & " addr1_buffer = "& Convert_SLV_To_Hex_String(addr1_buffer) & "outputs: " & " R_addr1_414_resized= "  & Convert_SLV_To_Hex_String(R_addr1_414_resized));
      --
    end process; 
    -- equivalence array_obj_ref_415_index_1_resize
    process(addr1_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr1_buffer;
      ov := iv(13 downto 0);
      R_addr1_414_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_415_root_address_inst flow-through 
    process(array_obj_ref_415_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_415_root_address_inst:flowthrough  inputs: " & " array_obj_ref_415_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_415_final_offset) & "outputs: " & " array_obj_ref_415_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_415_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_415_root_address_inst
    process(array_obj_ref_415_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_415_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_415_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_422_index_1_rename flow-through 
    process(R_addr2_421_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_422_index_1_rename:flowthrough  inputs: " & " R_addr2_421_resized = "& Convert_SLV_To_Hex_String(R_addr2_421_resized) & "outputs: " & " R_addr2_421_scaled= "  & Convert_SLV_To_Hex_String(R_addr2_421_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_422_index_1_rename
    process(R_addr2_421_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr2_421_resized;
      ov(13 downto 0) := iv;
      R_addr2_421_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_422_index_1_resize flow-through 
    process(R_addr2_421_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_422_index_1_resize:flowthrough  inputs: " & " addr2_buffer = "& Convert_SLV_To_Hex_String(addr2_buffer) & "outputs: " & " R_addr2_421_resized= "  & Convert_SLV_To_Hex_String(R_addr2_421_resized));
      --
    end process; 
    -- equivalence array_obj_ref_422_index_1_resize
    process(addr2_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr2_buffer;
      ov := iv(13 downto 0);
      R_addr2_421_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_422_root_address_inst flow-through 
    process(array_obj_ref_422_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_422_root_address_inst:flowthrough  inputs: " & " array_obj_ref_422_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_422_final_offset) & "outputs: " & " array_obj_ref_422_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_422_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_422_root_address_inst
    process(array_obj_ref_422_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_422_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_422_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_429_index_1_rename flow-through 
    process(R_addr3_428_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_429_index_1_rename:flowthrough  inputs: " & " R_addr3_428_resized = "& Convert_SLV_To_Hex_String(R_addr3_428_resized) & "outputs: " & " R_addr3_428_scaled= "  & Convert_SLV_To_Hex_String(R_addr3_428_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_429_index_1_rename
    process(R_addr3_428_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr3_428_resized;
      ov(13 downto 0) := iv;
      R_addr3_428_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_429_index_1_resize flow-through 
    process(R_addr3_428_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_429_index_1_resize:flowthrough  inputs: " & " addr3_buffer = "& Convert_SLV_To_Hex_String(addr3_buffer) & "outputs: " & " R_addr3_428_resized= "  & Convert_SLV_To_Hex_String(R_addr3_428_resized));
      --
    end process; 
    -- equivalence array_obj_ref_429_index_1_resize
    process(addr3_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr3_buffer;
      ov := iv(13 downto 0);
      R_addr3_428_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_429_root_address_inst flow-through 
    process(array_obj_ref_429_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_429_root_address_inst:flowthrough  inputs: " & " array_obj_ref_429_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_429_final_offset) & "outputs: " & " array_obj_ref_429_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_429_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_429_root_address_inst
    process(array_obj_ref_429_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_429_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_429_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_436_index_1_rename flow-through 
    process(R_addr4_435_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_436_index_1_rename:flowthrough  inputs: " & " R_addr4_435_resized = "& Convert_SLV_To_Hex_String(R_addr4_435_resized) & "outputs: " & " R_addr4_435_scaled= "  & Convert_SLV_To_Hex_String(R_addr4_435_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_436_index_1_rename
    process(R_addr4_435_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr4_435_resized;
      ov(13 downto 0) := iv;
      R_addr4_435_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_436_index_1_resize flow-through 
    process(R_addr4_435_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_436_index_1_resize:flowthrough  inputs: " & " addr4_buffer = "& Convert_SLV_To_Hex_String(addr4_buffer) & "outputs: " & " R_addr4_435_resized= "  & Convert_SLV_To_Hex_String(R_addr4_435_resized));
      --
    end process; 
    -- equivalence array_obj_ref_436_index_1_resize
    process(addr4_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr4_buffer;
      ov := iv(13 downto 0);
      R_addr4_435_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_436_root_address_inst flow-through 
    process(array_obj_ref_436_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_436_root_address_inst:flowthrough  inputs: " & " array_obj_ref_436_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_436_final_offset) & "outputs: " & " array_obj_ref_436_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_436_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_436_root_address_inst
    process(array_obj_ref_436_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_436_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_436_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1363_addr_0 flow-through 
    process(ptr_deref_1363_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1363_addr_0:flowthrough  inputs: " & " ptr_deref_1363_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1363_root_address) & "outputs: " & " ptr_deref_1363_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1363_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1363_addr_0
    process(ptr_deref_1363_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1363_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1363_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1363_base_resize flow-through 
    process(ptr_deref_1363_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1363_base_resize:flowthrough  inputs: " & " myptr5_1359_delayed_8_0_1361 = "& Convert_SLV_To_Hex_String(myptr5_1359_delayed_8_0_1361) & "outputs: " & " ptr_deref_1363_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1363_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1363_base_resize
    process(myptr5_1359_delayed_8_0_1361) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr5_1359_delayed_8_0_1361;
      ov := iv(13 downto 0);
      ptr_deref_1363_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1363_gather_scatter flow-through 
    process(ptr_deref_1363_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1363_gather_scatter:flowthrough  inputs: " & " CONCAT_u32_u64_1374_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_1374_wire) & "outputs: " & " ptr_deref_1363_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1363_data_0));
      --
    end process; 
    -- equivalence ptr_deref_1363_gather_scatter
    process(CONCAT_u32_u64_1374_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1374_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1363_data_0 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1363_root_address_inst flow-through 
    process(ptr_deref_1363_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1363_root_address_inst:flowthrough  inputs: " & " ptr_deref_1363_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1363_resized_base_address) & "outputs: " & " ptr_deref_1363_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1363_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1363_root_address_inst
    process(ptr_deref_1363_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1363_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1363_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1389_addr_0 flow-through 
    process(ptr_deref_1389_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1389_addr_0:flowthrough  inputs: " & " ptr_deref_1389_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1389_root_address) & "outputs: " & " ptr_deref_1389_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1389_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1389_addr_0
    process(ptr_deref_1389_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1389_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1389_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1389_base_resize flow-through 
    process(ptr_deref_1389_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1389_base_resize:flowthrough  inputs: " & " myptr6_1382_delayed_8_0_1387 = "& Convert_SLV_To_Hex_String(myptr6_1382_delayed_8_0_1387) & "outputs: " & " ptr_deref_1389_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1389_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1389_base_resize
    process(myptr6_1382_delayed_8_0_1387) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr6_1382_delayed_8_0_1387;
      ov := iv(13 downto 0);
      ptr_deref_1389_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1389_gather_scatter flow-through 
    process(ptr_deref_1389_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1389_gather_scatter:flowthrough  inputs: " & " CONCAT_u32_u64_1400_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_1400_wire) & "outputs: " & " ptr_deref_1389_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1389_data_0));
      --
    end process; 
    -- equivalence ptr_deref_1389_gather_scatter
    process(CONCAT_u32_u64_1400_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1400_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1389_data_0 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1389_root_address_inst flow-through 
    process(ptr_deref_1389_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1389_root_address_inst:flowthrough  inputs: " & " ptr_deref_1389_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1389_resized_base_address) & "outputs: " & " ptr_deref_1389_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1389_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1389_root_address_inst
    process(ptr_deref_1389_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1389_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1389_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1415_addr_0 flow-through 
    process(ptr_deref_1415_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1415_addr_0:flowthrough  inputs: " & " ptr_deref_1415_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1415_root_address) & "outputs: " & " ptr_deref_1415_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1415_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1415_addr_0
    process(ptr_deref_1415_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1415_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1415_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1415_base_resize flow-through 
    process(ptr_deref_1415_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1415_base_resize:flowthrough  inputs: " & " myptr7_1405_delayed_8_0_1413 = "& Convert_SLV_To_Hex_String(myptr7_1405_delayed_8_0_1413) & "outputs: " & " ptr_deref_1415_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1415_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1415_base_resize
    process(myptr7_1405_delayed_8_0_1413) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr7_1405_delayed_8_0_1413;
      ov := iv(13 downto 0);
      ptr_deref_1415_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1415_gather_scatter flow-through 
    process(ptr_deref_1415_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1415_gather_scatter:flowthrough  inputs: " & " CONCAT_u32_u64_1426_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_1426_wire) & "outputs: " & " ptr_deref_1415_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1415_data_0));
      --
    end process; 
    -- equivalence ptr_deref_1415_gather_scatter
    process(CONCAT_u32_u64_1426_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1426_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1415_data_0 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1415_root_address_inst flow-through 
    process(ptr_deref_1415_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1415_root_address_inst:flowthrough  inputs: " & " ptr_deref_1415_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1415_resized_base_address) & "outputs: " & " ptr_deref_1415_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1415_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1415_root_address_inst
    process(ptr_deref_1415_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1415_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1415_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1441_addr_0 flow-through 
    process(ptr_deref_1441_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1441_addr_0:flowthrough  inputs: " & " ptr_deref_1441_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1441_root_address) & "outputs: " & " ptr_deref_1441_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1441_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1441_addr_0
    process(ptr_deref_1441_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1441_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1441_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1441_base_resize flow-through 
    process(ptr_deref_1441_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1441_base_resize:flowthrough  inputs: " & " myptr8_1428_delayed_8_0_1439 = "& Convert_SLV_To_Hex_String(myptr8_1428_delayed_8_0_1439) & "outputs: " & " ptr_deref_1441_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1441_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1441_base_resize
    process(myptr8_1428_delayed_8_0_1439) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr8_1428_delayed_8_0_1439;
      ov := iv(13 downto 0);
      ptr_deref_1441_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1441_gather_scatter flow-through 
    process(ptr_deref_1441_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1441_gather_scatter:flowthrough  inputs: " & " CONCAT_u32_u64_1452_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_1452_wire) & "outputs: " & " ptr_deref_1441_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1441_data_0));
      --
    end process; 
    -- equivalence ptr_deref_1441_gather_scatter
    process(CONCAT_u32_u64_1452_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1452_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1441_data_0 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1441_root_address_inst flow-through 
    process(ptr_deref_1441_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1441_root_address_inst:flowthrough  inputs: " & " ptr_deref_1441_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1441_resized_base_address) & "outputs: " & " ptr_deref_1441_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1441_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1441_root_address_inst
    process(ptr_deref_1441_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1441_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1441_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_441_addr_0 flow-through 
    process(ptr_deref_441_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_441_addr_0:flowthrough  inputs: " & " ptr_deref_441_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_441_root_address) & "outputs: " & " ptr_deref_441_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_441_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_441_addr_0
    process(ptr_deref_441_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_441_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_441_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_441_base_resize flow-through 
    process(ptr_deref_441_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_441_base_resize:flowthrough  inputs: " & " myptr1_417 = "& Convert_SLV_To_Hex_String(myptr1_417) & "outputs: " & " ptr_deref_441_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_441_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_441_base_resize
    process(myptr1_417) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr1_417;
      ov := iv(13 downto 0);
      ptr_deref_441_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_441_gather_scatter flow-through 
    process(c1_442) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_441_gather_scatter:flowthrough  inputs: " & " ptr_deref_441_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_441_data_0) & "outputs: " & " c1_442= "  & Convert_SLV_To_Hex_String(c1_442));
      --
    end process; 
    -- equivalence ptr_deref_441_gather_scatter
    process(ptr_deref_441_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_441_data_0;
      ov(255 downto 0) := iv;
      c1_442 <= ov(255 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_441_root_address_inst flow-through 
    process(ptr_deref_441_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_441_root_address_inst:flowthrough  inputs: " & " ptr_deref_441_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_441_resized_base_address) & "outputs: " & " ptr_deref_441_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_441_root_address));
      --
    end process; 
    -- equivalence ptr_deref_441_root_address_inst
    process(ptr_deref_441_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_441_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_441_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_445_addr_0 flow-through 
    process(ptr_deref_445_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_445_addr_0:flowthrough  inputs: " & " ptr_deref_445_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_445_root_address) & "outputs: " & " ptr_deref_445_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_445_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_445_addr_0
    process(ptr_deref_445_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_445_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_445_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_445_base_resize flow-through 
    process(ptr_deref_445_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_445_base_resize:flowthrough  inputs: " & " myptr2_424 = "& Convert_SLV_To_Hex_String(myptr2_424) & "outputs: " & " ptr_deref_445_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_445_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_445_base_resize
    process(myptr2_424) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr2_424;
      ov := iv(13 downto 0);
      ptr_deref_445_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_445_gather_scatter flow-through 
    process(c2_446) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_445_gather_scatter:flowthrough  inputs: " & " ptr_deref_445_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_445_data_0) & "outputs: " & " c2_446= "  & Convert_SLV_To_Hex_String(c2_446));
      --
    end process; 
    -- equivalence ptr_deref_445_gather_scatter
    process(ptr_deref_445_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_445_data_0;
      ov(255 downto 0) := iv;
      c2_446 <= ov(255 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_445_root_address_inst flow-through 
    process(ptr_deref_445_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_445_root_address_inst:flowthrough  inputs: " & " ptr_deref_445_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_445_resized_base_address) & "outputs: " & " ptr_deref_445_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_445_root_address));
      --
    end process; 
    -- equivalence ptr_deref_445_root_address_inst
    process(ptr_deref_445_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_445_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_445_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_449_addr_0 flow-through 
    process(ptr_deref_449_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_449_addr_0:flowthrough  inputs: " & " ptr_deref_449_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_449_root_address) & "outputs: " & " ptr_deref_449_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_449_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_449_addr_0
    process(ptr_deref_449_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_449_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_449_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_449_base_resize flow-through 
    process(ptr_deref_449_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_449_base_resize:flowthrough  inputs: " & " myptr3_431 = "& Convert_SLV_To_Hex_String(myptr3_431) & "outputs: " & " ptr_deref_449_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_449_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_449_base_resize
    process(myptr3_431) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr3_431;
      ov := iv(13 downto 0);
      ptr_deref_449_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_449_gather_scatter flow-through 
    process(c3_450) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_449_gather_scatter:flowthrough  inputs: " & " ptr_deref_449_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_449_data_0) & "outputs: " & " c3_450= "  & Convert_SLV_To_Hex_String(c3_450));
      --
    end process; 
    -- equivalence ptr_deref_449_gather_scatter
    process(ptr_deref_449_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_449_data_0;
      ov(255 downto 0) := iv;
      c3_450 <= ov(255 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_449_root_address_inst flow-through 
    process(ptr_deref_449_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_449_root_address_inst:flowthrough  inputs: " & " ptr_deref_449_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_449_resized_base_address) & "outputs: " & " ptr_deref_449_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_449_root_address));
      --
    end process; 
    -- equivalence ptr_deref_449_root_address_inst
    process(ptr_deref_449_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_449_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_449_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_453_addr_0 flow-through 
    process(ptr_deref_453_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_453_addr_0:flowthrough  inputs: " & " ptr_deref_453_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_453_root_address) & "outputs: " & " ptr_deref_453_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_453_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_453_addr_0
    process(ptr_deref_453_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_453_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_453_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_453_base_resize flow-through 
    process(ptr_deref_453_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_453_base_resize:flowthrough  inputs: " & " myptr4_438 = "& Convert_SLV_To_Hex_String(myptr4_438) & "outputs: " & " ptr_deref_453_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_453_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_453_base_resize
    process(myptr4_438) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr4_438;
      ov := iv(13 downto 0);
      ptr_deref_453_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_453_gather_scatter flow-through 
    process(c4_454) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_453_gather_scatter:flowthrough  inputs: " & " ptr_deref_453_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_453_data_0) & "outputs: " & " c4_454= "  & Convert_SLV_To_Hex_String(c4_454));
      --
    end process; 
    -- equivalence ptr_deref_453_gather_scatter
    process(ptr_deref_453_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_453_data_0;
      ov(255 downto 0) := iv;
      c4_454 <= ov(255 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_453_root_address_inst flow-through 
    process(ptr_deref_453_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_453_root_address_inst:flowthrough  inputs: " & " ptr_deref_453_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_453_resized_base_address) & "outputs: " & " ptr_deref_453_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_453_root_address));
      --
    end process; 
    -- equivalence ptr_deref_453_root_address_inst
    process(ptr_deref_453_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_453_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_453_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for split-operator ADD_u32_u32_1381_inst flow-through 
    process(ADD_u32_u32_1381_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ADD_u32_u32_1381_inst:flowthrough inputs: " & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & " konst_1380_wire_constant = "& Convert_SLV_To_Hex_String(konst_1380_wire_constant) & " outputs:" & " ADD_u32_u32_1381_wire= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_1381_wire));
      --
    end process; 
    -- binary operator ADD_u32_u32_1381_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1380_wire_constant, tmp_var);
      ADD_u32_u32_1381_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1407_inst flow-through 
    process(ADD_u32_u32_1407_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ADD_u32_u32_1407_inst:flowthrough inputs: " & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & " konst_1406_wire_constant = "& Convert_SLV_To_Hex_String(konst_1406_wire_constant) & " outputs:" & " ADD_u32_u32_1407_wire= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_1407_wire));
      --
    end process; 
    -- binary operator ADD_u32_u32_1407_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1406_wire_constant, tmp_var);
      ADD_u32_u32_1407_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u32_u32_1433_inst flow-through 
    process(ADD_u32_u32_1433_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ADD_u32_u32_1433_inst:flowthrough inputs: " & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & " konst_1432_wire_constant = "& Convert_SLV_To_Hex_String(konst_1432_wire_constant) & " outputs:" & " ADD_u32_u32_1433_wire= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_1433_wire));
      --
    end process; 
    -- binary operator ADD_u32_u32_1433_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1432_wire_constant, tmp_var);
      ADD_u32_u32_1433_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_1368_inst flow-through 
    process(CONCAT_u16_u32_1368_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u16_u32_1368_inst:flowthrough inputs: " & " type_cast_1365_wire = "& Convert_SLV_To_Hex_String(type_cast_1365_wire) & " type_cast_1367_wire = "& Convert_SLV_To_Hex_String(type_cast_1367_wire) & " outputs:" & " CONCAT_u16_u32_1368_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_1368_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_1368_inst
    process(type_cast_1365_wire, type_cast_1367_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1365_wire, type_cast_1367_wire, tmp_var);
      CONCAT_u16_u32_1368_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_1373_inst flow-through 
    process(CONCAT_u16_u32_1373_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u16_u32_1373_inst:flowthrough inputs: " & " type_cast_1370_wire = "& Convert_SLV_To_Hex_String(type_cast_1370_wire) & " type_cast_1372_wire = "& Convert_SLV_To_Hex_String(type_cast_1372_wire) & " outputs:" & " CONCAT_u16_u32_1373_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_1373_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_1373_inst
    process(type_cast_1370_wire, type_cast_1372_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1370_wire, type_cast_1372_wire, tmp_var);
      CONCAT_u16_u32_1373_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_1394_inst flow-through 
    process(CONCAT_u16_u32_1394_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u16_u32_1394_inst:flowthrough inputs: " & " type_cast_1391_wire = "& Convert_SLV_To_Hex_String(type_cast_1391_wire) & " type_cast_1393_wire = "& Convert_SLV_To_Hex_String(type_cast_1393_wire) & " outputs:" & " CONCAT_u16_u32_1394_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_1394_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_1394_inst
    process(type_cast_1391_wire, type_cast_1393_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1391_wire, type_cast_1393_wire, tmp_var);
      CONCAT_u16_u32_1394_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_1399_inst flow-through 
    process(CONCAT_u16_u32_1399_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u16_u32_1399_inst:flowthrough inputs: " & " type_cast_1396_wire = "& Convert_SLV_To_Hex_String(type_cast_1396_wire) & " type_cast_1398_wire = "& Convert_SLV_To_Hex_String(type_cast_1398_wire) & " outputs:" & " CONCAT_u16_u32_1399_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_1399_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_1399_inst
    process(type_cast_1396_wire, type_cast_1398_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1396_wire, type_cast_1398_wire, tmp_var);
      CONCAT_u16_u32_1399_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_1420_inst flow-through 
    process(CONCAT_u16_u32_1420_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u16_u32_1420_inst:flowthrough inputs: " & " type_cast_1417_wire = "& Convert_SLV_To_Hex_String(type_cast_1417_wire) & " type_cast_1419_wire = "& Convert_SLV_To_Hex_String(type_cast_1419_wire) & " outputs:" & " CONCAT_u16_u32_1420_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_1420_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_1420_inst
    process(type_cast_1417_wire, type_cast_1419_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1417_wire, type_cast_1419_wire, tmp_var);
      CONCAT_u16_u32_1420_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_1425_inst flow-through 
    process(CONCAT_u16_u32_1425_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u16_u32_1425_inst:flowthrough inputs: " & " type_cast_1422_wire = "& Convert_SLV_To_Hex_String(type_cast_1422_wire) & " type_cast_1424_wire = "& Convert_SLV_To_Hex_String(type_cast_1424_wire) & " outputs:" & " CONCAT_u16_u32_1425_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_1425_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_1425_inst
    process(type_cast_1422_wire, type_cast_1424_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1422_wire, type_cast_1424_wire, tmp_var);
      CONCAT_u16_u32_1425_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_1446_inst flow-through 
    process(CONCAT_u16_u32_1446_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u16_u32_1446_inst:flowthrough inputs: " & " type_cast_1443_wire = "& Convert_SLV_To_Hex_String(type_cast_1443_wire) & " type_cast_1445_wire = "& Convert_SLV_To_Hex_String(type_cast_1445_wire) & " outputs:" & " CONCAT_u16_u32_1446_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_1446_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_1446_inst
    process(type_cast_1443_wire, type_cast_1445_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1443_wire, type_cast_1445_wire, tmp_var);
      CONCAT_u16_u32_1446_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_1451_inst flow-through 
    process(CONCAT_u16_u32_1451_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u16_u32_1451_inst:flowthrough inputs: " & " type_cast_1448_wire = "& Convert_SLV_To_Hex_String(type_cast_1448_wire) & " type_cast_1450_wire = "& Convert_SLV_To_Hex_String(type_cast_1450_wire) & " outputs:" & " CONCAT_u16_u32_1451_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_1451_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_1451_inst
    process(type_cast_1448_wire, type_cast_1450_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1448_wire, type_cast_1450_wire, tmp_var);
      CONCAT_u16_u32_1451_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u64_1374_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u32_u64_1374_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u32_u64_1374_inst:started:   inputs: " & " CONCAT_u16_u32_1368_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_1368_wire) & " CONCAT_u16_u32_1373_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_1373_wire));
          --
        end if; 
        if CONCAT_u32_u64_1374_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u32_u64_1374_inst:finished:  outputs: " & " CONCAT_u32_u64_1374_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_1374_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (11) : CONCAT_u32_u64_1374_inst 
    ApConcat_group_11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1368_wire & CONCAT_u16_u32_1373_wire;
      CONCAT_u32_u64_1374_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1374_inst_req_0;
      CONCAT_u32_u64_1374_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1374_inst_req_1;
      CONCAT_u32_u64_1374_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_11_gI: SplitGuardInterface generic map(name => "ApConcat_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- logger for split-operator CONCAT_u32_u64_1400_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u32_u64_1400_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u32_u64_1400_inst:started:   inputs: " & " CONCAT_u16_u32_1394_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_1394_wire) & " CONCAT_u16_u32_1399_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_1399_wire));
          --
        end if; 
        if CONCAT_u32_u64_1400_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u32_u64_1400_inst:finished:  outputs: " & " CONCAT_u32_u64_1400_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_1400_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (12) : CONCAT_u32_u64_1400_inst 
    ApConcat_group_12: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1394_wire & CONCAT_u16_u32_1399_wire;
      CONCAT_u32_u64_1400_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1400_inst_req_0;
      CONCAT_u32_u64_1400_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1400_inst_req_1;
      CONCAT_u32_u64_1400_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_12_gI: SplitGuardInterface generic map(name => "ApConcat_group_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- logger for split-operator CONCAT_u32_u64_1426_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u32_u64_1426_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u32_u64_1426_inst:started:   inputs: " & " CONCAT_u16_u32_1420_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_1420_wire) & " CONCAT_u16_u32_1425_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_1425_wire));
          --
        end if; 
        if CONCAT_u32_u64_1426_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u32_u64_1426_inst:finished:  outputs: " & " CONCAT_u32_u64_1426_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_1426_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (13) : CONCAT_u32_u64_1426_inst 
    ApConcat_group_13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1420_wire & CONCAT_u16_u32_1425_wire;
      CONCAT_u32_u64_1426_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1426_inst_req_0;
      CONCAT_u32_u64_1426_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1426_inst_req_1;
      CONCAT_u32_u64_1426_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_13_gI: SplitGuardInterface generic map(name => "ApConcat_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- logger for split-operator CONCAT_u32_u64_1452_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u32_u64_1452_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u32_u64_1452_inst:started:   inputs: " & " CONCAT_u16_u32_1446_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_1446_wire) & " CONCAT_u16_u32_1451_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_1451_wire));
          --
        end if; 
        if CONCAT_u32_u64_1452_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:CONCAT_u32_u64_1452_inst:finished:  outputs: " & " CONCAT_u32_u64_1452_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_1452_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (14) : CONCAT_u32_u64_1452_inst 
    ApConcat_group_14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1446_wire & CONCAT_u16_u32_1451_wire;
      CONCAT_u32_u64_1452_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1452_inst_req_0;
      CONCAT_u32_u64_1452_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1452_inst_req_1;
      CONCAT_u32_u64_1452_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_14_gI: SplitGuardInterface generic map(name => "ApConcat_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- logger for split-operator SGT_i16_u1_1003_inst flow-through 
    process(SGT_i16_u1_1003_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1003_inst:flowthrough inputs: " & " a32_847 = "& Convert_SLV_To_Hex_String(a32_847) & " a42_911 = "& Convert_SLV_To_Hex_String(a42_911) & " outputs:" & " SGT_i16_u1_1003_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1003_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1003_inst
    process(a32_847, a42_911) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a32_847, a42_911, tmp_var);
      SGT_i16_u1_1003_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1011_inst flow-through 
    process(SGT_i16_u1_1011_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1011_inst:flowthrough inputs: " & " t21_999 = "& Convert_SLV_To_Hex_String(t21_999) & " t22_1007 = "& Convert_SLV_To_Hex_String(t22_1007) & " outputs:" & " SGT_i16_u1_1011_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1011_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1011_inst
    process(t21_999, t22_1007) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t21_999, t22_1007, tmp_var);
      SGT_i16_u1_1011_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1019_inst flow-through 
    process(SGT_i16_u1_1019_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1019_inst:flowthrough inputs: " & " a13_723 = "& Convert_SLV_To_Hex_String(a13_723) & " a23_787 = "& Convert_SLV_To_Hex_String(a23_787) & " outputs:" & " SGT_i16_u1_1019_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1019_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1019_inst
    process(a13_723, a23_787) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a13_723, a23_787, tmp_var);
      SGT_i16_u1_1019_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1027_inst flow-through 
    process(SGT_i16_u1_1027_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1027_inst:flowthrough inputs: " & " a33_851 = "& Convert_SLV_To_Hex_String(a33_851) & " a43_915 = "& Convert_SLV_To_Hex_String(a43_915) & " outputs:" & " SGT_i16_u1_1027_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1027_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1027_inst
    process(a33_851, a43_915) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a33_851, a43_915, tmp_var);
      SGT_i16_u1_1027_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1035_inst flow-through 
    process(SGT_i16_u1_1035_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1035_inst:flowthrough inputs: " & " t31_1023 = "& Convert_SLV_To_Hex_String(t31_1023) & " t32_1031 = "& Convert_SLV_To_Hex_String(t32_1031) & " outputs:" & " SGT_i16_u1_1035_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1035_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1035_inst
    process(t31_1023, t32_1031) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t31_1023, t32_1031, tmp_var);
      SGT_i16_u1_1035_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1043_inst flow-through 
    process(SGT_i16_u1_1043_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1043_inst:flowthrough inputs: " & " a14_727 = "& Convert_SLV_To_Hex_String(a14_727) & " a24_791 = "& Convert_SLV_To_Hex_String(a24_791) & " outputs:" & " SGT_i16_u1_1043_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1043_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1043_inst
    process(a14_727, a24_791) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a14_727, a24_791, tmp_var);
      SGT_i16_u1_1043_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1051_inst flow-through 
    process(SGT_i16_u1_1051_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1051_inst:flowthrough inputs: " & " a34_855 = "& Convert_SLV_To_Hex_String(a34_855) & " a44_919 = "& Convert_SLV_To_Hex_String(a44_919) & " outputs:" & " SGT_i16_u1_1051_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1051_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1051_inst
    process(a34_855, a44_919) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a34_855, a44_919, tmp_var);
      SGT_i16_u1_1051_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1059_inst flow-through 
    process(SGT_i16_u1_1059_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1059_inst:flowthrough inputs: " & " t41_1047 = "& Convert_SLV_To_Hex_String(t41_1047) & " t42_1055 = "& Convert_SLV_To_Hex_String(t42_1055) & " outputs:" & " SGT_i16_u1_1059_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1059_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1059_inst
    process(t41_1047, t42_1055) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t41_1047, t42_1055, tmp_var);
      SGT_i16_u1_1059_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1067_inst flow-through 
    process(SGT_i16_u1_1067_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1067_inst:flowthrough inputs: " & " a15_731 = "& Convert_SLV_To_Hex_String(a15_731) & " a25_795 = "& Convert_SLV_To_Hex_String(a25_795) & " outputs:" & " SGT_i16_u1_1067_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1067_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1067_inst
    process(a15_731, a25_795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a15_731, a25_795, tmp_var);
      SGT_i16_u1_1067_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1075_inst flow-through 
    process(SGT_i16_u1_1075_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1075_inst:flowthrough inputs: " & " a35_859 = "& Convert_SLV_To_Hex_String(a35_859) & " a45_923 = "& Convert_SLV_To_Hex_String(a45_923) & " outputs:" & " SGT_i16_u1_1075_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1075_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1075_inst
    process(a35_859, a45_923) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a35_859, a45_923, tmp_var);
      SGT_i16_u1_1075_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1083_inst flow-through 
    process(SGT_i16_u1_1083_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1083_inst:flowthrough inputs: " & " t51_1071 = "& Convert_SLV_To_Hex_String(t51_1071) & " t52_1079 = "& Convert_SLV_To_Hex_String(t52_1079) & " outputs:" & " SGT_i16_u1_1083_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1083_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1083_inst
    process(t51_1071, t52_1079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t51_1071, t52_1079, tmp_var);
      SGT_i16_u1_1083_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1091_inst flow-through 
    process(SGT_i16_u1_1091_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1091_inst:flowthrough inputs: " & " a16_735 = "& Convert_SLV_To_Hex_String(a16_735) & " a26_799 = "& Convert_SLV_To_Hex_String(a26_799) & " outputs:" & " SGT_i16_u1_1091_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1091_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1091_inst
    process(a16_735, a26_799) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a16_735, a26_799, tmp_var);
      SGT_i16_u1_1091_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1099_inst flow-through 
    process(SGT_i16_u1_1099_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1099_inst:flowthrough inputs: " & " a36_863 = "& Convert_SLV_To_Hex_String(a36_863) & " a46_927 = "& Convert_SLV_To_Hex_String(a46_927) & " outputs:" & " SGT_i16_u1_1099_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1099_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1099_inst
    process(a36_863, a46_927) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a36_863, a46_927, tmp_var);
      SGT_i16_u1_1099_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1107_inst flow-through 
    process(SGT_i16_u1_1107_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1107_inst:flowthrough inputs: " & " t61_1095 = "& Convert_SLV_To_Hex_String(t61_1095) & " t62_1103 = "& Convert_SLV_To_Hex_String(t62_1103) & " outputs:" & " SGT_i16_u1_1107_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1107_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1107_inst
    process(t61_1095, t62_1103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t61_1095, t62_1103, tmp_var);
      SGT_i16_u1_1107_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1115_inst flow-through 
    process(SGT_i16_u1_1115_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1115_inst:flowthrough inputs: " & " a17_739 = "& Convert_SLV_To_Hex_String(a17_739) & " a27_803 = "& Convert_SLV_To_Hex_String(a27_803) & " outputs:" & " SGT_i16_u1_1115_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1115_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1115_inst
    process(a17_739, a27_803) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a17_739, a27_803, tmp_var);
      SGT_i16_u1_1115_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1123_inst flow-through 
    process(SGT_i16_u1_1123_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1123_inst:flowthrough inputs: " & " a37_867 = "& Convert_SLV_To_Hex_String(a37_867) & " a47_931 = "& Convert_SLV_To_Hex_String(a47_931) & " outputs:" & " SGT_i16_u1_1123_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1123_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1123_inst
    process(a37_867, a47_931) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a37_867, a47_931, tmp_var);
      SGT_i16_u1_1123_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1131_inst flow-through 
    process(SGT_i16_u1_1131_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1131_inst:flowthrough inputs: " & " t71_1119 = "& Convert_SLV_To_Hex_String(t71_1119) & " t72_1127 = "& Convert_SLV_To_Hex_String(t72_1127) & " outputs:" & " SGT_i16_u1_1131_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1131_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1131_inst
    process(t71_1119, t72_1127) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t71_1119, t72_1127, tmp_var);
      SGT_i16_u1_1131_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1139_inst flow-through 
    process(SGT_i16_u1_1139_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1139_inst:flowthrough inputs: " & " a18_743 = "& Convert_SLV_To_Hex_String(a18_743) & " a28_807 = "& Convert_SLV_To_Hex_String(a28_807) & " outputs:" & " SGT_i16_u1_1139_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1139_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1139_inst
    process(a18_743, a28_807) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a18_743, a28_807, tmp_var);
      SGT_i16_u1_1139_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1147_inst flow-through 
    process(SGT_i16_u1_1147_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1147_inst:flowthrough inputs: " & " a38_871 = "& Convert_SLV_To_Hex_String(a38_871) & " a48_935 = "& Convert_SLV_To_Hex_String(a48_935) & " outputs:" & " SGT_i16_u1_1147_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1147_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1147_inst
    process(a38_871, a48_935) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a38_871, a48_935, tmp_var);
      SGT_i16_u1_1147_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1155_inst flow-through 
    process(SGT_i16_u1_1155_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1155_inst:flowthrough inputs: " & " t81_1143 = "& Convert_SLV_To_Hex_String(t81_1143) & " t82_1151 = "& Convert_SLV_To_Hex_String(t82_1151) & " outputs:" & " SGT_i16_u1_1155_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1155_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1155_inst
    process(t81_1143, t82_1151) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t81_1143, t82_1151, tmp_var);
      SGT_i16_u1_1155_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1163_inst flow-through 
    process(SGT_i16_u1_1163_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1163_inst:flowthrough inputs: " & " a19_747 = "& Convert_SLV_To_Hex_String(a19_747) & " a29_811 = "& Convert_SLV_To_Hex_String(a29_811) & " outputs:" & " SGT_i16_u1_1163_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1163_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1163_inst
    process(a19_747, a29_811) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a19_747, a29_811, tmp_var);
      SGT_i16_u1_1163_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1171_inst flow-through 
    process(SGT_i16_u1_1171_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1171_inst:flowthrough inputs: " & " a39_875 = "& Convert_SLV_To_Hex_String(a39_875) & " a49_939 = "& Convert_SLV_To_Hex_String(a49_939) & " outputs:" & " SGT_i16_u1_1171_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1171_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1171_inst
    process(a39_875, a49_939) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a39_875, a49_939, tmp_var);
      SGT_i16_u1_1171_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1179_inst flow-through 
    process(SGT_i16_u1_1179_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1179_inst:flowthrough inputs: " & " t91_1167 = "& Convert_SLV_To_Hex_String(t91_1167) & " t92_1175 = "& Convert_SLV_To_Hex_String(t92_1175) & " outputs:" & " SGT_i16_u1_1179_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1179_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1179_inst
    process(t91_1167, t92_1175) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t91_1167, t92_1175, tmp_var);
      SGT_i16_u1_1179_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1187_inst flow-through 
    process(SGT_i16_u1_1187_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1187_inst:flowthrough inputs: " & " a110_751 = "& Convert_SLV_To_Hex_String(a110_751) & " a210_815 = "& Convert_SLV_To_Hex_String(a210_815) & " outputs:" & " SGT_i16_u1_1187_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1187_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1187_inst
    process(a110_751, a210_815) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a110_751, a210_815, tmp_var);
      SGT_i16_u1_1187_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1195_inst flow-through 
    process(SGT_i16_u1_1195_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1195_inst:flowthrough inputs: " & " a310_879 = "& Convert_SLV_To_Hex_String(a310_879) & " a410_943 = "& Convert_SLV_To_Hex_String(a410_943) & " outputs:" & " SGT_i16_u1_1195_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1195_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1195_inst
    process(a310_879, a410_943) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a310_879, a410_943, tmp_var);
      SGT_i16_u1_1195_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1203_inst flow-through 
    process(SGT_i16_u1_1203_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1203_inst:flowthrough inputs: " & " t101_1191 = "& Convert_SLV_To_Hex_String(t101_1191) & " t102_1199 = "& Convert_SLV_To_Hex_String(t102_1199) & " outputs:" & " SGT_i16_u1_1203_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1203_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1203_inst
    process(t101_1191, t102_1199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t101_1191, t102_1199, tmp_var);
      SGT_i16_u1_1203_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1211_inst flow-through 
    process(SGT_i16_u1_1211_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1211_inst:flowthrough inputs: " & " a111_755 = "& Convert_SLV_To_Hex_String(a111_755) & " a211_819 = "& Convert_SLV_To_Hex_String(a211_819) & " outputs:" & " SGT_i16_u1_1211_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1211_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1211_inst
    process(a111_755, a211_819) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a111_755, a211_819, tmp_var);
      SGT_i16_u1_1211_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1219_inst flow-through 
    process(SGT_i16_u1_1219_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1219_inst:flowthrough inputs: " & " a311_883 = "& Convert_SLV_To_Hex_String(a311_883) & " a411_947 = "& Convert_SLV_To_Hex_String(a411_947) & " outputs:" & " SGT_i16_u1_1219_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1219_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1219_inst
    process(a311_883, a411_947) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a311_883, a411_947, tmp_var);
      SGT_i16_u1_1219_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1227_inst flow-through 
    process(SGT_i16_u1_1227_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1227_inst:flowthrough inputs: " & " t111_1215 = "& Convert_SLV_To_Hex_String(t111_1215) & " t112_1223 = "& Convert_SLV_To_Hex_String(t112_1223) & " outputs:" & " SGT_i16_u1_1227_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1227_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1227_inst
    process(t111_1215, t112_1223) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t111_1215, t112_1223, tmp_var);
      SGT_i16_u1_1227_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1235_inst flow-through 
    process(SGT_i16_u1_1235_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1235_inst:flowthrough inputs: " & " a112_759 = "& Convert_SLV_To_Hex_String(a112_759) & " a212_823 = "& Convert_SLV_To_Hex_String(a212_823) & " outputs:" & " SGT_i16_u1_1235_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1235_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1235_inst
    process(a112_759, a212_823) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a112_759, a212_823, tmp_var);
      SGT_i16_u1_1235_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1243_inst flow-through 
    process(SGT_i16_u1_1243_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1243_inst:flowthrough inputs: " & " a312_887 = "& Convert_SLV_To_Hex_String(a312_887) & " a412_951 = "& Convert_SLV_To_Hex_String(a412_951) & " outputs:" & " SGT_i16_u1_1243_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1243_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1243_inst
    process(a312_887, a412_951) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a312_887, a412_951, tmp_var);
      SGT_i16_u1_1243_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1251_inst flow-through 
    process(SGT_i16_u1_1251_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1251_inst:flowthrough inputs: " & " t121_1239 = "& Convert_SLV_To_Hex_String(t121_1239) & " t122_1247 = "& Convert_SLV_To_Hex_String(t122_1247) & " outputs:" & " SGT_i16_u1_1251_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1251_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1251_inst
    process(t121_1239, t122_1247) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t121_1239, t122_1247, tmp_var);
      SGT_i16_u1_1251_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1259_inst flow-through 
    process(SGT_i16_u1_1259_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1259_inst:flowthrough inputs: " & " a113_763 = "& Convert_SLV_To_Hex_String(a113_763) & " a213_827 = "& Convert_SLV_To_Hex_String(a213_827) & " outputs:" & " SGT_i16_u1_1259_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1259_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1259_inst
    process(a113_763, a213_827) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a113_763, a213_827, tmp_var);
      SGT_i16_u1_1259_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1267_inst flow-through 
    process(SGT_i16_u1_1267_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1267_inst:flowthrough inputs: " & " a313_891 = "& Convert_SLV_To_Hex_String(a313_891) & " a413_955 = "& Convert_SLV_To_Hex_String(a413_955) & " outputs:" & " SGT_i16_u1_1267_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1267_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1267_inst
    process(a313_891, a413_955) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a313_891, a413_955, tmp_var);
      SGT_i16_u1_1267_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1275_inst flow-through 
    process(SGT_i16_u1_1275_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1275_inst:flowthrough inputs: " & " t131_1263 = "& Convert_SLV_To_Hex_String(t131_1263) & " t132_1271 = "& Convert_SLV_To_Hex_String(t132_1271) & " outputs:" & " SGT_i16_u1_1275_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1275_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1275_inst
    process(t131_1263, t132_1271) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t131_1263, t132_1271, tmp_var);
      SGT_i16_u1_1275_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1283_inst flow-through 
    process(SGT_i16_u1_1283_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1283_inst:flowthrough inputs: " & " a114_767 = "& Convert_SLV_To_Hex_String(a114_767) & " a214_831 = "& Convert_SLV_To_Hex_String(a214_831) & " outputs:" & " SGT_i16_u1_1283_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1283_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1283_inst
    process(a114_767, a214_831) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a114_767, a214_831, tmp_var);
      SGT_i16_u1_1283_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1291_inst flow-through 
    process(SGT_i16_u1_1291_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1291_inst:flowthrough inputs: " & " a314_895 = "& Convert_SLV_To_Hex_String(a314_895) & " a414_959 = "& Convert_SLV_To_Hex_String(a414_959) & " outputs:" & " SGT_i16_u1_1291_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1291_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1291_inst
    process(a314_895, a414_959) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a314_895, a414_959, tmp_var);
      SGT_i16_u1_1291_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1299_inst flow-through 
    process(SGT_i16_u1_1299_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1299_inst:flowthrough inputs: " & " t141_1287 = "& Convert_SLV_To_Hex_String(t141_1287) & " t142_1295 = "& Convert_SLV_To_Hex_String(t142_1295) & " outputs:" & " SGT_i16_u1_1299_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1299_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1299_inst
    process(t141_1287, t142_1295) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t141_1287, t142_1295, tmp_var);
      SGT_i16_u1_1299_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1307_inst flow-through 
    process(SGT_i16_u1_1307_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1307_inst:flowthrough inputs: " & " a115_771 = "& Convert_SLV_To_Hex_String(a115_771) & " a215_835 = "& Convert_SLV_To_Hex_String(a215_835) & " outputs:" & " SGT_i16_u1_1307_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1307_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1307_inst
    process(a115_771, a215_835) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a115_771, a215_835, tmp_var);
      SGT_i16_u1_1307_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1315_inst flow-through 
    process(SGT_i16_u1_1315_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1315_inst:flowthrough inputs: " & " a315_899 = "& Convert_SLV_To_Hex_String(a315_899) & " a415_963 = "& Convert_SLV_To_Hex_String(a415_963) & " outputs:" & " SGT_i16_u1_1315_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1315_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1315_inst
    process(a315_899, a415_963) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a315_899, a415_963, tmp_var);
      SGT_i16_u1_1315_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1323_inst flow-through 
    process(SGT_i16_u1_1323_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1323_inst:flowthrough inputs: " & " t151_1311 = "& Convert_SLV_To_Hex_String(t151_1311) & " t152_1319 = "& Convert_SLV_To_Hex_String(t152_1319) & " outputs:" & " SGT_i16_u1_1323_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1323_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1323_inst
    process(t151_1311, t152_1319) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t151_1311, t152_1319, tmp_var);
      SGT_i16_u1_1323_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1331_inst flow-through 
    process(SGT_i16_u1_1331_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1331_inst:flowthrough inputs: " & " a116_775 = "& Convert_SLV_To_Hex_String(a116_775) & " a216_839 = "& Convert_SLV_To_Hex_String(a216_839) & " outputs:" & " SGT_i16_u1_1331_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1331_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1331_inst
    process(a116_775, a216_839) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a116_775, a216_839, tmp_var);
      SGT_i16_u1_1331_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1339_inst flow-through 
    process(SGT_i16_u1_1339_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1339_inst:flowthrough inputs: " & " a316_903 = "& Convert_SLV_To_Hex_String(a316_903) & " a416_967 = "& Convert_SLV_To_Hex_String(a416_967) & " outputs:" & " SGT_i16_u1_1339_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1339_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1339_inst
    process(a316_903, a416_967) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a316_903, a416_967, tmp_var);
      SGT_i16_u1_1339_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_1347_inst flow-through 
    process(SGT_i16_u1_1347_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_1347_inst:flowthrough inputs: " & " t161_1335 = "& Convert_SLV_To_Hex_String(t161_1335) & " t162_1343 = "& Convert_SLV_To_Hex_String(t162_1343) & " outputs:" & " SGT_i16_u1_1347_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_1347_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_1347_inst
    process(t161_1335, t162_1343) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t161_1335, t162_1343, tmp_var);
      SGT_i16_u1_1347_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_971_inst flow-through 
    process(SGT_i16_u1_971_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_971_inst:flowthrough inputs: " & " a11_715 = "& Convert_SLV_To_Hex_String(a11_715) & " a21_779 = "& Convert_SLV_To_Hex_String(a21_779) & " outputs:" & " SGT_i16_u1_971_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_971_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_971_inst
    process(a11_715, a21_779) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a11_715, a21_779, tmp_var);
      SGT_i16_u1_971_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_979_inst flow-through 
    process(SGT_i16_u1_979_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_979_inst:flowthrough inputs: " & " a31_843 = "& Convert_SLV_To_Hex_String(a31_843) & " a41_907 = "& Convert_SLV_To_Hex_String(a41_907) & " outputs:" & " SGT_i16_u1_979_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_979_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_979_inst
    process(a31_843, a41_907) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a31_843, a41_907, tmp_var);
      SGT_i16_u1_979_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_987_inst flow-through 
    process(SGT_i16_u1_987_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_987_inst:flowthrough inputs: " & " t11_975 = "& Convert_SLV_To_Hex_String(t11_975) & " t12_983 = "& Convert_SLV_To_Hex_String(t12_983) & " outputs:" & " SGT_i16_u1_987_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_987_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_987_inst
    process(t11_975, t12_983) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t11_975, t12_983, tmp_var);
      SGT_i16_u1_987_wire <= tmp_var; --
    end process;
    -- logger for split-operator SGT_i16_u1_995_inst flow-through 
    process(SGT_i16_u1_995_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:SGT_i16_u1_995_inst:flowthrough inputs: " & " a12_719 = "& Convert_SLV_To_Hex_String(a12_719) & " a22_783 = "& Convert_SLV_To_Hex_String(a22_783) & " outputs:" & " SGT_i16_u1_995_wire= "  & Convert_SLV_To_Hex_String(SGT_i16_u1_995_wire));
      --
    end process; 
    -- binary operator SGT_i16_u1_995_inst
    process(a12_719, a22_783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a12_719, a22_783, tmp_var);
      SGT_i16_u1_995_wire <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_1356_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1356_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1356_index_offset:started:   inputs: " & " R_addr_1355_scaled = "& Convert_SLV_To_Hex_String(R_addr_1355_scaled) & " array_obj_ref_1356_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1356_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1356_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1356_index_offset:finished:  outputs: " & " array_obj_ref_1356_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1356_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (63) : array_obj_ref_1356_index_offset 
    ApIntAdd_group_63: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_1355_scaled;
      array_obj_ref_1356_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1356_index_offset_req_0;
      array_obj_ref_1356_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1356_index_offset_req_1;
      array_obj_ref_1356_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_63_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_63_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_63",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- logger for split-operator array_obj_ref_1382_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1382_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1382_index_offset:started:   inputs: " & " ADD_u32_u32_1381_scaled = "& Convert_SLV_To_Hex_String(ADD_u32_u32_1381_scaled) & " array_obj_ref_1382_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1382_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1382_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1382_index_offset:finished:  outputs: " & " array_obj_ref_1382_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1382_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (64) : array_obj_ref_1382_index_offset 
    ApIntAdd_group_64: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1381_scaled;
      array_obj_ref_1382_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1382_index_offset_req_0;
      array_obj_ref_1382_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1382_index_offset_req_1;
      array_obj_ref_1382_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_64_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_64_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_64",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- logger for split-operator array_obj_ref_1408_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1408_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1408_index_offset:started:   inputs: " & " ADD_u32_u32_1407_scaled = "& Convert_SLV_To_Hex_String(ADD_u32_u32_1407_scaled) & " array_obj_ref_1408_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1408_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1408_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1408_index_offset:finished:  outputs: " & " array_obj_ref_1408_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1408_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (65) : array_obj_ref_1408_index_offset 
    ApIntAdd_group_65: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1407_scaled;
      array_obj_ref_1408_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1408_index_offset_req_0;
      array_obj_ref_1408_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1408_index_offset_req_1;
      array_obj_ref_1408_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_65_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_65_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_65",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- logger for split-operator array_obj_ref_1434_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1434_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1434_index_offset:started:   inputs: " & " ADD_u32_u32_1433_scaled = "& Convert_SLV_To_Hex_String(ADD_u32_u32_1433_scaled) & " array_obj_ref_1434_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1434_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1434_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_1434_index_offset:finished:  outputs: " & " array_obj_ref_1434_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1434_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (66) : array_obj_ref_1434_index_offset 
    ApIntAdd_group_66: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1433_scaled;
      array_obj_ref_1434_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1434_index_offset_req_0;
      array_obj_ref_1434_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1434_index_offset_req_1;
      array_obj_ref_1434_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_66_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_66_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_66",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- logger for split-operator array_obj_ref_415_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_415_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_415_index_offset:started:   inputs: " & " R_addr1_414_scaled = "& Convert_SLV_To_Hex_String(R_addr1_414_scaled) & " array_obj_ref_415_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_415_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_415_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_415_index_offset:finished:  outputs: " & " array_obj_ref_415_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_415_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (67) : array_obj_ref_415_index_offset 
    ApIntAdd_group_67: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr1_414_scaled;
      array_obj_ref_415_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_415_index_offset_req_0;
      array_obj_ref_415_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_415_index_offset_req_1;
      array_obj_ref_415_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_67_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_67_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_67",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- logger for split-operator array_obj_ref_422_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_422_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_422_index_offset:started:   inputs: " & " R_addr2_421_scaled = "& Convert_SLV_To_Hex_String(R_addr2_421_scaled) & " array_obj_ref_422_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_422_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_422_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_422_index_offset:finished:  outputs: " & " array_obj_ref_422_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_422_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (68) : array_obj_ref_422_index_offset 
    ApIntAdd_group_68: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr2_421_scaled;
      array_obj_ref_422_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_422_index_offset_req_0;
      array_obj_ref_422_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_422_index_offset_req_1;
      array_obj_ref_422_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_68_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_68_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_68",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- logger for split-operator array_obj_ref_429_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_429_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_429_index_offset:started:   inputs: " & " R_addr3_428_scaled = "& Convert_SLV_To_Hex_String(R_addr3_428_scaled) & " array_obj_ref_429_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_429_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_429_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_429_index_offset:finished:  outputs: " & " array_obj_ref_429_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_429_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (69) : array_obj_ref_429_index_offset 
    ApIntAdd_group_69: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr3_428_scaled;
      array_obj_ref_429_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_429_index_offset_req_0;
      array_obj_ref_429_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_429_index_offset_req_1;
      array_obj_ref_429_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_69_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_69_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_69",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- logger for split-operator array_obj_ref_436_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_436_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_436_index_offset:started:   inputs: " & " R_addr4_435_scaled = "& Convert_SLV_To_Hex_String(R_addr4_435_scaled) & " array_obj_ref_436_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_436_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_436_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:array_obj_ref_436_index_offset:finished:  outputs: " & " array_obj_ref_436_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_436_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (70) : array_obj_ref_436_index_offset 
    ApIntAdd_group_70: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr4_435_scaled;
      array_obj_ref_436_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_436_index_offset_req_0;
      array_obj_ref_436_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_436_index_offset_req_1;
      array_obj_ref_436_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_70_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_70_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_70",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- logger for split-operator ptr_deref_449_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_449_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_449_load_0:started:   inputs: " & " ptr_deref_449_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_449_word_address_0));
          --
        end if; 
        if ptr_deref_449_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_449_load_0:finished:  outputs: " & " ptr_deref_449_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_449_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_445_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_445_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_445_load_0:started:   inputs: " & " ptr_deref_445_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_445_word_address_0));
          --
        end if; 
        if ptr_deref_445_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_445_load_0:finished:  outputs: " & " ptr_deref_445_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_445_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_453_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_453_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_453_load_0:started:   inputs: " & " ptr_deref_453_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_453_word_address_0));
          --
        end if; 
        if ptr_deref_453_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_453_load_0:finished:  outputs: " & " ptr_deref_453_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_453_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_441_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_441_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_441_load_0:started:   inputs: " & " ptr_deref_441_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_441_word_address_0));
          --
        end if; 
        if ptr_deref_441_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_441_load_0:finished:  outputs: " & " ptr_deref_441_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_441_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : ptr_deref_449_load_0 ptr_deref_445_load_0 ptr_deref_453_load_0 ptr_deref_441_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(1023 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_449_load_0_req_0,
        ptr_deref_449_load_0_ack_0,
        ptr_deref_449_load_0_req_1,
        ptr_deref_449_load_0_ack_1,
        "ptr_deref_449_load_0",
        "memory_space_1" ,
        ptr_deref_449_data_0,
        ptr_deref_449_word_address_0,
        "ptr_deref_449_data_0",
        "ptr_deref_449_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_445_load_0_req_0,
        ptr_deref_445_load_0_ack_0,
        ptr_deref_445_load_0_req_1,
        ptr_deref_445_load_0_ack_1,
        "ptr_deref_445_load_0",
        "memory_space_1" ,
        ptr_deref_445_data_0,
        ptr_deref_445_word_address_0,
        "ptr_deref_445_data_0",
        "ptr_deref_445_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_453_load_0_req_0,
        ptr_deref_453_load_0_ack_0,
        ptr_deref_453_load_0_req_1,
        ptr_deref_453_load_0_ack_1,
        "ptr_deref_453_load_0",
        "memory_space_1" ,
        ptr_deref_453_data_0,
        ptr_deref_453_word_address_0,
        "ptr_deref_453_data_0",
        "ptr_deref_453_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_441_load_0_req_0,
        ptr_deref_441_load_0_ack_0,
        ptr_deref_441_load_0_req_1,
        ptr_deref_441_load_0_ack_1,
        "ptr_deref_441_load_0",
        "memory_space_1" ,
        ptr_deref_441_data_0,
        ptr_deref_441_word_address_0,
        "ptr_deref_441_data_0",
        "ptr_deref_441_word_address_0" -- 
      );
      reqL_unguarded(3) <= ptr_deref_449_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_445_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_453_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_441_load_0_req_0;
      ptr_deref_449_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_445_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_453_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_441_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_449_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_445_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_453_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_441_load_0_req_1;
      ptr_deref_449_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_445_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_453_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_441_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_449_word_address_0 & ptr_deref_445_word_address_0 & ptr_deref_453_word_address_0 & ptr_deref_441_word_address_0;
      ptr_deref_449_data_0 <= data_out(1023 downto 768);
      ptr_deref_445_data_0 <= data_out(767 downto 512);
      ptr_deref_453_data_0 <= data_out(511 downto 256);
      ptr_deref_441_data_0 <= data_out(255 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 256,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(255 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator ptr_deref_1363_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1363_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1363_store_0:started:   inputs: " & " ptr_deref_1363_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1363_word_address_0) & " ptr_deref_1363_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1363_data_0));
          --
        end if; 
        if ptr_deref_1363_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1363_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_1415_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1415_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1415_store_0:started:   inputs: " & " ptr_deref_1415_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1415_word_address_0) & " ptr_deref_1415_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1415_data_0));
          --
        end if; 
        if ptr_deref_1415_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1415_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_1389_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1389_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1389_store_0:started:   inputs: " & " ptr_deref_1389_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1389_word_address_0) & " ptr_deref_1389_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1389_data_0));
          --
        end if; 
        if ptr_deref_1389_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1389_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_1441_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1441_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1441_store_0:started:   inputs: " & " ptr_deref_1441_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1441_word_address_0) & " ptr_deref_1441_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1441_data_0));
          --
        end if; 
        if ptr_deref_1441_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:maxPool4:DP:ptr_deref_1441_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1363_store_0_req_0,
      ptr_deref_1363_store_0_ack_0,
      ptr_deref_1363_store_0_req_1,
      ptr_deref_1363_store_0_ack_1,
      "ptr_deref_1363_store_0",
      "memory_space_0" ,
      ptr_deref_1363_data_0,
      ptr_deref_1363_word_address_0,
      "ptr_deref_1363_data_0",
      "ptr_deref_1363_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1415_store_0_req_0,
      ptr_deref_1415_store_0_ack_0,
      ptr_deref_1415_store_0_req_1,
      ptr_deref_1415_store_0_ack_1,
      "ptr_deref_1415_store_0",
      "memory_space_0" ,
      ptr_deref_1415_data_0,
      ptr_deref_1415_word_address_0,
      "ptr_deref_1415_data_0",
      "ptr_deref_1415_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1389_store_0_req_0,
      ptr_deref_1389_store_0_ack_0,
      ptr_deref_1389_store_0_req_1,
      ptr_deref_1389_store_0_ack_1,
      "ptr_deref_1389_store_0",
      "memory_space_0" ,
      ptr_deref_1389_data_0,
      ptr_deref_1389_word_address_0,
      "ptr_deref_1389_data_0",
      "ptr_deref_1389_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1441_store_0_req_0,
      ptr_deref_1441_store_0_ack_0,
      ptr_deref_1441_store_0_req_1,
      ptr_deref_1441_store_0_ack_1,
      "ptr_deref_1441_store_0",
      "memory_space_0" ,
      ptr_deref_1441_data_0,
      ptr_deref_1441_word_address_0,
      "ptr_deref_1441_data_0",
      "ptr_deref_1441_word_address_0" -- 
    );
    -- shared store operator group (0) : ptr_deref_1363_store_0 ptr_deref_1415_store_0 ptr_deref_1389_store_0 ptr_deref_1441_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(55 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 15, 2 => 15, 1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_1363_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1415_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1389_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1441_store_0_req_0;
      ptr_deref_1363_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1415_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1389_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1441_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_1363_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1415_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1389_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1441_store_0_req_1;
      ptr_deref_1363_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1415_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1389_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1441_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1363_word_address_0 & ptr_deref_1415_word_address_0 & ptr_deref_1389_word_address_0 & ptr_deref_1441_word_address_0;
      data_in <= ptr_deref_1363_data_0 & ptr_deref_1415_data_0 & ptr_deref_1389_data_0 & ptr_deref_1441_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 4,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end maxPool4_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendB;
architecture sendB_arch of sendB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendB_CP_3659_start: Boolean;
  signal sendB_CP_3659_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_1477_branch_ack_0 : boolean;
  signal ptr_deref_1469_load_0_req_0 : boolean;
  signal type_cast_1498_inst_ack_1 : boolean;
  signal ptr_deref_1469_load_0_req_1 : boolean;
  signal ptr_deref_1469_load_0_ack_1 : boolean;
  signal ptr_deref_1469_load_0_ack_0 : boolean;
  signal type_cast_1498_inst_req_0 : boolean;
  signal type_cast_1498_inst_ack_0 : boolean;
  signal type_cast_1498_inst_req_1 : boolean;
  signal if_stmt_1477_branch_ack_1 : boolean;
  signal if_stmt_1477_branch_req_0 : boolean;
  signal array_obj_ref_1534_index_offset_req_0 : boolean;
  signal array_obj_ref_1534_index_offset_ack_0 : boolean;
  signal array_obj_ref_1534_index_offset_req_1 : boolean;
  signal array_obj_ref_1534_index_offset_ack_1 : boolean;
  signal addr_of_1535_final_reg_req_0 : boolean;
  signal addr_of_1535_final_reg_ack_0 : boolean;
  signal addr_of_1535_final_reg_req_1 : boolean;
  signal addr_of_1535_final_reg_ack_1 : boolean;
  signal ptr_deref_1539_load_0_req_0 : boolean;
  signal ptr_deref_1539_load_0_ack_0 : boolean;
  signal ptr_deref_1539_load_0_req_1 : boolean;
  signal ptr_deref_1539_load_0_ack_1 : boolean;
  signal if_stmt_1557_branch_req_0 : boolean;
  signal if_stmt_1557_branch_ack_1 : boolean;
  signal if_stmt_1557_branch_ack_0 : boolean;
  signal if_stmt_1583_branch_req_0 : boolean;
  signal if_stmt_1583_branch_ack_1 : boolean;
  signal if_stmt_1583_branch_ack_0 : boolean;
  signal type_cast_1598_inst_req_0 : boolean;
  signal type_cast_1598_inst_ack_0 : boolean;
  signal type_cast_1598_inst_req_1 : boolean;
  signal type_cast_1598_inst_ack_1 : boolean;
  signal array_obj_ref_1633_index_offset_req_0 : boolean;
  signal array_obj_ref_1633_index_offset_ack_0 : boolean;
  signal array_obj_ref_1633_index_offset_req_1 : boolean;
  signal array_obj_ref_1633_index_offset_ack_1 : boolean;
  signal addr_of_1634_final_reg_req_0 : boolean;
  signal addr_of_1634_final_reg_ack_0 : boolean;
  signal addr_of_1634_final_reg_req_1 : boolean;
  signal addr_of_1634_final_reg_ack_1 : boolean;
  signal ptr_deref_1638_load_0_req_0 : boolean;
  signal ptr_deref_1638_load_0_ack_0 : boolean;
  signal ptr_deref_1638_load_0_req_1 : boolean;
  signal ptr_deref_1638_load_0_ack_1 : boolean;
  signal type_cast_1642_inst_req_0 : boolean;
  signal type_cast_1642_inst_ack_0 : boolean;
  signal type_cast_1642_inst_req_1 : boolean;
  signal type_cast_1642_inst_ack_1 : boolean;
  signal type_cast_1652_inst_req_0 : boolean;
  signal type_cast_1652_inst_ack_0 : boolean;
  signal type_cast_1652_inst_req_1 : boolean;
  signal type_cast_1652_inst_ack_1 : boolean;
  signal type_cast_1662_inst_req_0 : boolean;
  signal type_cast_1662_inst_ack_0 : boolean;
  signal type_cast_1662_inst_req_1 : boolean;
  signal type_cast_1662_inst_ack_1 : boolean;
  signal type_cast_1672_inst_req_0 : boolean;
  signal type_cast_1672_inst_ack_0 : boolean;
  signal type_cast_1672_inst_req_1 : boolean;
  signal type_cast_1672_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1677_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1677_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1677_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1677_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1680_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1680_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1680_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1680_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1683_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1683_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1683_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1683_inst_ack_1 : boolean;
  signal if_stmt_1697_branch_req_0 : boolean;
  signal if_stmt_1697_branch_ack_1 : boolean;
  signal if_stmt_1697_branch_ack_0 : boolean;
  signal phi_stmt_1515_req_0 : boolean;
  signal phi_stmt_1522_req_0 : boolean;
  signal type_cast_1521_inst_req_0 : boolean;
  signal type_cast_1521_inst_ack_0 : boolean;
  signal type_cast_1521_inst_req_1 : boolean;
  signal type_cast_1521_inst_ack_1 : boolean;
  signal phi_stmt_1515_req_1 : boolean;
  signal type_cast_1528_inst_req_0 : boolean;
  signal type_cast_1528_inst_ack_0 : boolean;
  signal type_cast_1528_inst_req_1 : boolean;
  signal type_cast_1528_inst_ack_1 : boolean;
  signal phi_stmt_1522_req_1 : boolean;
  signal phi_stmt_1515_ack_0 : boolean;
  signal phi_stmt_1522_ack_0 : boolean;
  signal type_cast_1567_inst_req_0 : boolean;
  signal type_cast_1567_inst_ack_0 : boolean;
  signal type_cast_1567_inst_req_1 : boolean;
  signal type_cast_1567_inst_ack_1 : boolean;
  signal phi_stmt_1564_req_0 : boolean;
  signal type_cast_1571_inst_req_0 : boolean;
  signal type_cast_1571_inst_ack_0 : boolean;
  signal type_cast_1571_inst_req_1 : boolean;
  signal type_cast_1571_inst_ack_1 : boolean;
  signal phi_stmt_1568_req_0 : boolean;
  signal type_cast_1575_inst_req_0 : boolean;
  signal type_cast_1575_inst_ack_0 : boolean;
  signal type_cast_1575_inst_req_1 : boolean;
  signal type_cast_1575_inst_ack_1 : boolean;
  signal phi_stmt_1572_req_0 : boolean;
  signal phi_stmt_1564_ack_0 : boolean;
  signal phi_stmt_1568_ack_0 : boolean;
  signal phi_stmt_1572_ack_0 : boolean;
  signal phi_stmt_1621_req_0 : boolean;
  signal type_cast_1627_inst_req_0 : boolean;
  signal type_cast_1627_inst_ack_0 : boolean;
  signal type_cast_1627_inst_req_1 : boolean;
  signal type_cast_1627_inst_ack_1 : boolean;
  signal phi_stmt_1621_req_1 : boolean;
  signal phi_stmt_1621_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendB_CP_3659_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_3659_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendB_CP_3659_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_3659_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,sendB_CP_3659_start,"sendB cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,sendB_CP_3659_symbol, "sendB cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendB_CP_3659: Block -- control-path 
    signal sendB_CP_3659_elements: BooleanArray(83 downto 0);
    -- 
  begin -- 
    sendB_CP_3659_elements(0) <= sendB_CP_3659_start;
    sendB_CP_3659_symbol <= sendB_CP_3659_elements(83);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (31) 
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1460/$entry
      -- CP-element group 0: 	 branch_block_stmt_1460/branch_block_stmt_1460__entry__
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476__entry__
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/$entry
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_word_addrgen/root_register_req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1469_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1469_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_3738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(0), ack => ptr_deref_1469_load_0_req_0); -- 
    cr_3749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(0), ack => ptr_deref_1469_load_0_req_1); -- 
    -- CP-element group 1:  merge  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	76 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	17 
    -- CP-element group 1: 	18 
    -- CP-element group 1:  members (13) 
      -- CP-element group 1: 	 branch_block_stmt_1460/R_cmp1357_1584_place
      -- CP-element group 1: 	 branch_block_stmt_1460/merge_stmt_1563__exit__
      -- CP-element group 1: 	 branch_block_stmt_1460/assign_stmt_1582__entry__
      -- CP-element group 1: 	 branch_block_stmt_1460/assign_stmt_1582__exit__
      -- CP-element group 1: 	 branch_block_stmt_1460/if_stmt_1583__entry__
      -- CP-element group 1: 	 branch_block_stmt_1460/assign_stmt_1582/$entry
      -- CP-element group 1: 	 branch_block_stmt_1460/assign_stmt_1582/$exit
      -- CP-element group 1: 	 branch_block_stmt_1460/if_stmt_1583_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1460/if_stmt_1583_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_1460/if_stmt_1583_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_1460/if_stmt_1583_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_1460/if_stmt_1583_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1460/if_stmt_1583_else_link/$entry
      -- 
    -- logger for CP element group sendB_CP_3659_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1583_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_3920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(1), ack => if_stmt_1583_branch_req_0); -- 
    sendB_CP_3659_elements(1) <= sendB_CP_3659_elements(76);
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Sample/word_access_start/$exit
      -- CP-element group 2: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Sample/word_access_start/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Sample/word_access_start/word_0/ra
      -- CP-element group 2: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_sample_completed_
      -- 
    -- logger for CP element group sendB_CP_3659_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1469_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1469_load_0_ack_0, ack => sendB_CP_3659_elements(2)); -- 
    -- CP-element group 3:  branch  transition  place  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	5 
    -- CP-element group 3:  members (19) 
      -- CP-element group 3: 	 branch_block_stmt_1460/R_cmp60_1478_place
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/ptr_deref_1469_Merge/$entry
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/word_access_complete/word_0/ca
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/ptr_deref_1469_Merge/merge_ack
      -- CP-element group 3: 	 branch_block_stmt_1460/if_stmt_1477_dead_link/$entry
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/ptr_deref_1469_Merge/merge_req
      -- CP-element group 3: 	 branch_block_stmt_1460/if_stmt_1477_eval_test/$entry
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/word_access_complete/$exit
      -- CP-element group 3: 	 branch_block_stmt_1460/if_stmt_1477_eval_test/$exit
      -- CP-element group 3: 	 branch_block_stmt_1460/if_stmt_1477_eval_test/branch_req
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/ptr_deref_1469_Merge/$exit
      -- CP-element group 3: 	 branch_block_stmt_1460/if_stmt_1477_if_link/$entry
      -- CP-element group 3: 	 branch_block_stmt_1460/if_stmt_1477_else_link/$entry
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_Update/word_access_complete/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476__exit__
      -- CP-element group 3: 	 branch_block_stmt_1460/if_stmt_1477__entry__
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/$exit
      -- CP-element group 3: 	 branch_block_stmt_1460/assign_stmt_1466_to_assign_stmt_1476/ptr_deref_1469_update_completed_
      -- 
    -- logger for CP element group sendB_CP_3659_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1469_load_0_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1477_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_3750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1469_load_0_ack_1, ack => sendB_CP_3659_elements(3)); -- 
    branch_req_3763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(3), ack => if_stmt_1477_branch_req_0); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	83 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 branch_block_stmt_1460/entry_forx_xend54
      -- CP-element group 4: 	 branch_block_stmt_1460/if_stmt_1477_if_link/$exit
      -- CP-element group 4: 	 branch_block_stmt_1460/if_stmt_1477_if_link/if_choice_transition
      -- CP-element group 4: 	 branch_block_stmt_1460/entry_forx_xend54_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1460/entry_forx_xend54_PhiReq/$exit
      -- 
    -- logger for CP element group sendB_CP_3659_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1477_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_3768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1477_branch_ack_1, ack => sendB_CP_3659_elements(4)); -- 
    -- CP-element group 5:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	3 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (18) 
      -- CP-element group 5: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1460/if_stmt_1477_else_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1460/if_stmt_1477_else_link/else_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_1460/entry_bbx_xnph63
      -- CP-element group 5: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/$entry
      -- CP-element group 5: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1460/merge_stmt_1483__exit__
      -- CP-element group 5: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512__entry__
      -- CP-element group 5: 	 branch_block_stmt_1460/entry_bbx_xnph63_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1460/entry_bbx_xnph63_PhiReq/$exit
      -- CP-element group 5: 	 branch_block_stmt_1460/merge_stmt_1483_PhiReqMerge
      -- CP-element group 5: 	 branch_block_stmt_1460/merge_stmt_1483_PhiAck/$entry
      -- CP-element group 5: 	 branch_block_stmt_1460/merge_stmt_1483_PhiAck/$exit
      -- CP-element group 5: 	 branch_block_stmt_1460/merge_stmt_1483_PhiAck/dummy
      -- 
    -- logger for CP element group sendB_CP_3659_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1477_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1498_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1498_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_3772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1477_branch_ack_0, ack => sendB_CP_3659_elements(5)); -- 
    rr_3785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(5), ack => type_cast_1498_inst_req_0); -- 
    cr_3790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(5), ack => type_cast_1498_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1498_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1498_inst_ack_0, ack => sendB_CP_3659_elements(6)); -- 
    -- CP-element group 7:  fork  transition  place  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	49 
    -- CP-element group 7: 	50 
    -- CP-element group 7:  members (11) 
      -- CP-element group 7: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/$exit
      -- CP-element group 7: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512/type_cast_1498_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1460/assign_stmt_1489_to_assign_stmt_1512__exit__
      -- CP-element group 7: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody
      -- CP-element group 7: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/$entry
      -- CP-element group 7: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1515/$entry
      -- CP-element group 7: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1522/$entry
      -- CP-element group 7: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/$entry
      -- 
    -- logger for CP element group sendB_CP_3659_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1498_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1498_inst_ack_1, ack => sendB_CP_3659_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	62 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_final_index_sum_regn_sample_complete
      -- CP-element group 8: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_final_index_sum_regn_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:array_obj_ref_1534_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1534_index_offset_ack_0, ack => sendB_CP_3659_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	62 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (11) 
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_offset_calculated
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_final_index_sum_regn_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_final_index_sum_regn_Update/ack
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_base_plus_offset/$entry
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_base_plus_offset/$exit
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_base_plus_offset/sum_rename_req
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_base_plus_offset/sum_rename_ack
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_request/$entry
      -- CP-element group 9: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_request/req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:array_obj_ref_1534_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:addr_of_1535_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1534_index_offset_ack_1, ack => sendB_CP_3659_elements(9)); -- 
    req_3834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(9), ack => addr_of_1535_final_reg_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_request/$exit
      -- CP-element group 10: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_request/ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:addr_of_1535_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1535_final_reg_ack_0, ack => sendB_CP_3659_elements(10)); -- 
    -- CP-element group 11:  join  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	62 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (24) 
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_complete/$exit
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_complete/ack
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_base_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_base_address_resized
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_base_addr_resize/$entry
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_base_addr_resize/$exit
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_base_addr_resize/base_resize_req
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_base_addr_resize/base_resize_ack
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_base_plus_offset/$entry
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_base_plus_offset/$exit
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_base_plus_offset/sum_rename_req
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_base_plus_offset/sum_rename_ack
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_word_addrgen/$entry
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_word_addrgen/$exit
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_word_addrgen/root_register_req
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_word_addrgen/root_register_ack
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Sample/word_access_start/$entry
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Sample/word_access_start/word_0/$entry
      -- CP-element group 11: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group sendB_CP_3659_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:addr_of_1535_final_reg_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1539_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1535_final_reg_ack_1, ack => sendB_CP_3659_elements(11)); -- 
    rr_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(11), ack => ptr_deref_1539_load_0_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Sample/word_access_start/$exit
      -- CP-element group 12: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1539_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1539_load_0_ack_0, ack => sendB_CP_3659_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	62 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/word_access_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/ptr_deref_1539_Merge/$entry
      -- CP-element group 13: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/ptr_deref_1539_Merge/$exit
      -- CP-element group 13: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/ptr_deref_1539_Merge/merge_req
      -- CP-element group 13: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/ptr_deref_1539_Merge/merge_ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1539_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1539_load_0_ack_1, ack => sendB_CP_3659_elements(13)); -- 
    -- CP-element group 14:  branch  join  transition  place  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (10) 
      -- CP-element group 14: 	 branch_block_stmt_1460/R_exitcond_1558_place
      -- CP-element group 14: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/$exit
      -- CP-element group 14: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556__exit__
      -- CP-element group 14: 	 branch_block_stmt_1460/if_stmt_1557__entry__
      -- CP-element group 14: 	 branch_block_stmt_1460/if_stmt_1557_dead_link/$entry
      -- CP-element group 14: 	 branch_block_stmt_1460/if_stmt_1557_eval_test/$entry
      -- CP-element group 14: 	 branch_block_stmt_1460/if_stmt_1557_eval_test/$exit
      -- CP-element group 14: 	 branch_block_stmt_1460/if_stmt_1557_eval_test/branch_req
      -- CP-element group 14: 	 branch_block_stmt_1460/if_stmt_1557_if_link/$entry
      -- CP-element group 14: 	 branch_block_stmt_1460/if_stmt_1557_else_link/$entry
      -- 
    -- logger for CP element group sendB_CP_3659_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1557_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_3898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(14), ack => if_stmt_1557_branch_req_0); -- 
    sendB_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(8) & sendB_CP_3659_elements(13);
      gj_sendB_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	63 
    -- CP-element group 15: 	64 
    -- CP-element group 15: 	66 
    -- CP-element group 15: 	67 
    -- CP-element group 15: 	69 
    -- CP-element group 15: 	70 
    -- CP-element group 15:  members (28) 
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend
      -- CP-element group 15: 	 branch_block_stmt_1460/if_stmt_1557_if_link/$exit
      -- CP-element group 15: 	 branch_block_stmt_1460/if_stmt_1557_if_link/if_choice_transition
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/SplitProtocol/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/SplitProtocol/Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/SplitProtocol/Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/SplitProtocol/Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/SplitProtocol/Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/SplitProtocol/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/SplitProtocol/Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/SplitProtocol/Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/SplitProtocol/Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/SplitProtocol/Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/SplitProtocol/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/SplitProtocol/Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/SplitProtocol/Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/SplitProtocol/Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group sendB_CP_3659_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1557_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1567_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1567_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1571_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1571_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1575_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1575_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_3903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1557_branch_ack_1, ack => sendB_CP_3659_elements(15)); -- 
    rr_4287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(15), ack => type_cast_1567_inst_req_0); -- 
    cr_4292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(15), ack => type_cast_1567_inst_req_1); -- 
    rr_4310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(15), ack => type_cast_1571_inst_req_0); -- 
    cr_4315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(15), ack => type_cast_1571_inst_req_1); -- 
    rr_4333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(15), ack => type_cast_1575_inst_req_0); -- 
    cr_4338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(15), ack => type_cast_1575_inst_req_1); -- 
    -- CP-element group 16:  fork  transition  place  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	52 
    -- CP-element group 16: 	53 
    -- CP-element group 16: 	55 
    -- CP-element group 16: 	56 
    -- CP-element group 16:  members (20) 
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody
      -- CP-element group 16: 	 branch_block_stmt_1460/if_stmt_1557_else_link/$exit
      -- CP-element group 16: 	 branch_block_stmt_1460/if_stmt_1557_else_link/else_choice_transition
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group sendB_CP_3659_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1557_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1521_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1521_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1528_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1528_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_3907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1557_branch_ack_0, ack => sendB_CP_3659_elements(16)); -- 
    rr_4228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(16), ack => type_cast_1521_inst_req_0); -- 
    cr_4233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(16), ack => type_cast_1521_inst_req_1); -- 
    rr_4251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(16), ack => type_cast_1528_inst_req_0); -- 
    cr_4256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(16), ack => type_cast_1528_inst_req_1); -- 
    -- CP-element group 17:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	20 
    -- CP-element group 17:  members (18) 
      -- CP-element group 17: 	 branch_block_stmt_1460/forx_xend_bbx_xnph
      -- CP-element group 17: 	 branch_block_stmt_1460/merge_stmt_1589__exit__
      -- CP-element group 17: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618__entry__
      -- CP-element group 17: 	 branch_block_stmt_1460/if_stmt_1583_if_link/$exit
      -- CP-element group 17: 	 branch_block_stmt_1460/if_stmt_1583_if_link/if_choice_transition
      -- CP-element group 17: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/$entry
      -- CP-element group 17: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1460/forx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 17: 	 branch_block_stmt_1460/forx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 17: 	 branch_block_stmt_1460/merge_stmt_1589_PhiReqMerge
      -- CP-element group 17: 	 branch_block_stmt_1460/merge_stmt_1589_PhiAck/$entry
      -- CP-element group 17: 	 branch_block_stmt_1460/merge_stmt_1589_PhiAck/$exit
      -- CP-element group 17: 	 branch_block_stmt_1460/merge_stmt_1589_PhiAck/dummy
      -- 
    -- logger for CP element group sendB_CP_3659_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1583_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1598_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1598_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_3925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1583_branch_ack_1, ack => sendB_CP_3659_elements(17)); -- 
    rr_3942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(17), ack => type_cast_1598_inst_req_0); -- 
    cr_3947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(17), ack => type_cast_1598_inst_req_1); -- 
    -- CP-element group 18:  transition  place  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	83 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 branch_block_stmt_1460/forx_xend_forx_xend54
      -- CP-element group 18: 	 branch_block_stmt_1460/if_stmt_1583_else_link/$exit
      -- CP-element group 18: 	 branch_block_stmt_1460/if_stmt_1583_else_link/else_choice_transition
      -- CP-element group 18: 	 branch_block_stmt_1460/forx_xend_forx_xend54_PhiReq/$entry
      -- CP-element group 18: 	 branch_block_stmt_1460/forx_xend_forx_xend54_PhiReq/$exit
      -- 
    -- logger for CP element group sendB_CP_3659_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1583_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1583_branch_ack_0, ack => sendB_CP_3659_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1598_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1598_inst_ack_0, ack => sendB_CP_3659_elements(19)); -- 
    -- CP-element group 20:  transition  place  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	77 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618__exit__
      -- CP-element group 20: 	 branch_block_stmt_1460/bbx_xnph_forx_xbody15
      -- CP-element group 20: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/$exit
      -- CP-element group 20: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1460/assign_stmt_1594_to_assign_stmt_1618/type_cast_1598_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1460/bbx_xnph_forx_xbody15_PhiReq/$entry
      -- CP-element group 20: 	 branch_block_stmt_1460/bbx_xnph_forx_xbody15_PhiReq/phi_stmt_1621/$entry
      -- CP-element group 20: 	 branch_block_stmt_1460/bbx_xnph_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$entry
      -- 
    -- logger for CP element group sendB_CP_3659_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1598_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1598_inst_ack_1, ack => sendB_CP_3659_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	82 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	46 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_final_index_sum_regn_sample_complete
      -- CP-element group 21: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_final_index_sum_regn_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:array_obj_ref_1633_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1633_index_offset_ack_0, ack => sendB_CP_3659_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	82 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (11) 
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_root_address_calculated
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_offset_calculated
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_final_index_sum_regn_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_final_index_sum_regn_Update/ack
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_base_plus_offset/$entry
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_base_plus_offset/$exit
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_base_plus_offset/sum_rename_req
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_base_plus_offset/sum_rename_ack
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_request/$entry
      -- CP-element group 22: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_request/req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:array_obj_ref_1633_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:addr_of_1634_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1633_index_offset_ack_1, ack => sendB_CP_3659_elements(22)); -- 
    req_3991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(22), ack => addr_of_1634_final_reg_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_request/$exit
      -- CP-element group 23: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_request/ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:addr_of_1634_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1634_final_reg_ack_0, ack => sendB_CP_3659_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	82 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (24) 
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_complete/ack
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_base_address_calculated
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_word_address_calculated
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_root_address_calculated
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_base_address_resized
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_base_addr_resize/$entry
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_base_addr_resize/$exit
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_base_addr_resize/base_resize_req
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_base_addr_resize/base_resize_ack
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_base_plus_offset/$entry
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_base_plus_offset/$exit
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_base_plus_offset/sum_rename_req
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_base_plus_offset/sum_rename_ack
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_word_addrgen/$entry
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_word_addrgen/$exit
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_word_addrgen/root_register_req
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_word_addrgen/root_register_ack
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Sample/word_access_start/$entry
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Sample/word_access_start/word_0/$entry
      -- CP-element group 24: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group sendB_CP_3659_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:addr_of_1634_final_reg_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1638_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1634_final_reg_ack_1, ack => sendB_CP_3659_elements(24)); -- 
    rr_4030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(24), ack => ptr_deref_1638_load_0_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1638_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1638_load_0_ack_0, ack => sendB_CP_3659_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	82 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26: 	31 
    -- CP-element group 26: 	33 
    -- CP-element group 26:  members (21) 
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/ptr_deref_1638_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/ptr_deref_1638_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/ptr_deref_1638_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/ptr_deref_1638_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_Sample/rr
      -- 
    -- logger for CP element group sendB_CP_3659_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1638_load_0_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1642_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1652_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1662_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1672_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_4042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1638_load_0_ack_1, ack => sendB_CP_3659_elements(26)); -- 
    rr_4055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(26), ack => type_cast_1642_inst_req_0); -- 
    rr_4069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(26), ack => type_cast_1652_inst_req_0); -- 
    rr_4083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(26), ack => type_cast_1662_inst_req_0); -- 
    rr_4097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(26), ack => type_cast_1672_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1642_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1642_inst_ack_0, ack => sendB_CP_3659_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	82 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	43 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_Update/ca
      -- 
    -- logger for CP element group sendB_CP_3659_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1642_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1642_inst_ack_1, ack => sendB_CP_3659_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1652_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1652_inst_ack_0, ack => sendB_CP_3659_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	82 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	40 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_Update/ca
      -- 
    -- logger for CP element group sendB_CP_3659_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1652_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1652_inst_ack_1, ack => sendB_CP_3659_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1662_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1662_inst_ack_0, ack => sendB_CP_3659_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	82 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	37 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_Update/ca
      -- 
    -- logger for CP element group sendB_CP_3659_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1662_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1662_inst_ack_1, ack => sendB_CP_3659_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	26 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1672_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1672_inst_ack_0, ack => sendB_CP_3659_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	82 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_Sample/req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1672_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1674_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_4103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1672_inst_ack_1, ack => sendB_CP_3659_elements(34)); -- 
    req_4111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(34), ack => WPIPE_maxpool_output_pipe_1674_inst_req_0); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_Sample/ack
      -- CP-element group 35: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_Update/req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1674_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1674_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1674_inst_ack_0, ack => sendB_CP_3659_elements(35)); -- 
    req_4116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(35), ack => WPIPE_maxpool_output_pipe_1674_inst_req_1); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1674_Update/ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1674_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1674_inst_ack_1, ack => sendB_CP_3659_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	32 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_Sample/req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1677_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_4125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(37), ack => WPIPE_maxpool_output_pipe_1677_inst_req_0); -- 
    sendB_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(32) & sendB_CP_3659_elements(36);
      gj_sendB_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_Update/req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1677_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1677_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1677_inst_ack_0, ack => sendB_CP_3659_elements(38)); -- 
    req_4130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(38), ack => WPIPE_maxpool_output_pipe_1677_inst_req_1); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1677_Update/ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1677_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1677_inst_ack_1, ack => sendB_CP_3659_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	30 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_Sample/req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1680_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_4139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(40), ack => WPIPE_maxpool_output_pipe_1680_inst_req_0); -- 
    sendB_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(30) & sendB_CP_3659_elements(39);
      gj_sendB_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_Sample/ack
      -- CP-element group 41: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_Update/req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1680_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1680_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1680_inst_ack_0, ack => sendB_CP_3659_elements(41)); -- 
    req_4144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(41), ack => WPIPE_maxpool_output_pipe_1680_inst_req_1); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1680_Update/ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1680_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1680_inst_ack_1, ack => sendB_CP_3659_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	28 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_Sample/req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1683_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_4153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(43), ack => WPIPE_maxpool_output_pipe_1683_inst_req_0); -- 
    sendB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(28) & sendB_CP_3659_elements(42);
      gj_sendB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_update_start_
      -- CP-element group 44: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_Sample/ack
      -- CP-element group 44: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_Update/req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1683_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1683_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1683_inst_ack_0, ack => sendB_CP_3659_elements(44)); -- 
    req_4158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(44), ack => WPIPE_maxpool_output_pipe_1683_inst_req_1); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/WPIPE_maxpool_output_pipe_1683_Update/ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:WPIPE_maxpool_output_pipe_1683_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1683_inst_ack_1, ack => sendB_CP_3659_elements(45)); -- 
    -- CP-element group 46:  branch  join  transition  place  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	21 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (10) 
      -- CP-element group 46: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696__exit__
      -- CP-element group 46: 	 branch_block_stmt_1460/if_stmt_1697__entry__
      -- CP-element group 46: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/$exit
      -- CP-element group 46: 	 branch_block_stmt_1460/if_stmt_1697_dead_link/$entry
      -- CP-element group 46: 	 branch_block_stmt_1460/if_stmt_1697_eval_test/$entry
      -- CP-element group 46: 	 branch_block_stmt_1460/if_stmt_1697_eval_test/$exit
      -- CP-element group 46: 	 branch_block_stmt_1460/if_stmt_1697_eval_test/branch_req
      -- CP-element group 46: 	 branch_block_stmt_1460/R_exitcond7_1698_place
      -- CP-element group 46: 	 branch_block_stmt_1460/if_stmt_1697_if_link/$entry
      -- CP-element group 46: 	 branch_block_stmt_1460/if_stmt_1697_else_link/$entry
      -- 
    -- logger for CP element group sendB_CP_3659_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1697_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_4167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(46), ack => if_stmt_1697_branch_req_0); -- 
    sendB_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(21) & sendB_CP_3659_elements(45);
      gj_sendB_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  merge  transition  place  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	83 
    -- CP-element group 47:  members (13) 
      -- CP-element group 47: 	 branch_block_stmt_1460/merge_stmt_1703__exit__
      -- CP-element group 47: 	 branch_block_stmt_1460/forx_xend54x_xloopexit_forx_xend54
      -- CP-element group 47: 	 branch_block_stmt_1460/if_stmt_1697_if_link/$exit
      -- CP-element group 47: 	 branch_block_stmt_1460/if_stmt_1697_if_link/if_choice_transition
      -- CP-element group 47: 	 branch_block_stmt_1460/forx_xbody15_forx_xend54x_xloopexit
      -- CP-element group 47: 	 branch_block_stmt_1460/forx_xbody15_forx_xend54x_xloopexit_PhiReq/$entry
      -- CP-element group 47: 	 branch_block_stmt_1460/forx_xbody15_forx_xend54x_xloopexit_PhiReq/$exit
      -- CP-element group 47: 	 branch_block_stmt_1460/merge_stmt_1703_PhiReqMerge
      -- CP-element group 47: 	 branch_block_stmt_1460/merge_stmt_1703_PhiAck/$entry
      -- CP-element group 47: 	 branch_block_stmt_1460/merge_stmt_1703_PhiAck/$exit
      -- CP-element group 47: 	 branch_block_stmt_1460/merge_stmt_1703_PhiAck/dummy
      -- CP-element group 47: 	 branch_block_stmt_1460/forx_xend54x_xloopexit_forx_xend54_PhiReq/$entry
      -- CP-element group 47: 	 branch_block_stmt_1460/forx_xend54x_xloopexit_forx_xend54_PhiReq/$exit
      -- 
    -- logger for CP element group sendB_CP_3659_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1697_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_4172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1697_branch_ack_1, ack => sendB_CP_3659_elements(47)); -- 
    -- CP-element group 48:  fork  transition  place  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	78 
    -- CP-element group 48: 	79 
    -- CP-element group 48:  members (12) 
      -- CP-element group 48: 	 branch_block_stmt_1460/if_stmt_1697_else_link/$exit
      -- CP-element group 48: 	 branch_block_stmt_1460/if_stmt_1697_else_link/else_choice_transition
      -- CP-element group 48: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15
      -- CP-element group 48: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/$entry
      -- CP-element group 48: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/$entry
      -- CP-element group 48: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$entry
      -- CP-element group 48: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/$entry
      -- CP-element group 48: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/$entry
      -- CP-element group 48: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/rr
      -- CP-element group 48: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group sendB_CP_3659_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:if_stmt_1697_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1627_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1627_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_4176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1697_branch_ack_0, ack => sendB_CP_3659_elements(48)); -- 
    rr_4389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(48), ack => type_cast_1627_inst_req_0); -- 
    cr_4394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(48), ack => type_cast_1627_inst_req_1); -- 
    -- CP-element group 49:  transition  output  delay-element  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	7 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1515/$exit
      -- CP-element group 49: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$exit
      -- CP-element group 49: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1519_konst_delay_trans
      -- CP-element group 49: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1515_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1515_req_4201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1515_req_4201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(49), ack => phi_stmt_1515_req_0); -- 
    -- Element group sendB_CP_3659_elements(49) is a control-delay.
    cp_element_49_delay: control_delay_element  generic map(name => " 49_delay", delay_value => 1)  port map(req => sendB_CP_3659_elements(7), ack => sendB_CP_3659_elements(49), clk => clk, reset =>reset);
    -- CP-element group 50:  transition  output  delay-element  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	7 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1522/$exit
      -- CP-element group 50: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/$exit
      -- CP-element group 50: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1526_konst_delay_trans
      -- CP-element group 50: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1522_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1522_req_4209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1522_req_4209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(50), ack => phi_stmt_1522_req_0); -- 
    -- Element group sendB_CP_3659_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => sendB_CP_3659_elements(7), ack => sendB_CP_3659_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  transition  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1460/bbx_xnph63_forx_xbody_PhiReq/$exit
      -- 
    -- logger for CP element group sendB_CP_3659_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    sendB_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(49) & sendB_CP_3659_elements(50);
      gj_sendB_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	16 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (2) 
      -- CP-element group 52: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1521_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_0, ack => sendB_CP_3659_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	16 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group sendB_CP_3659_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1521_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_1, ack => sendB_CP_3659_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	58 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/$exit
      -- CP-element group 54: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$exit
      -- CP-element group 54: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/$exit
      -- CP-element group 54: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/$exit
      -- CP-element group 54: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1515/phi_stmt_1515_req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1515_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1515_req_4235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1515_req_4235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(54), ack => phi_stmt_1515_req_1); -- 
    sendB_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(52) & sendB_CP_3659_elements(53);
      gj_sendB_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	16 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1528_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1528_inst_ack_0, ack => sendB_CP_3659_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	16 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group sendB_CP_3659_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1528_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1528_inst_ack_1, ack => sendB_CP_3659_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/$exit
      -- CP-element group 57: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/$exit
      -- CP-element group 57: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/$exit
      -- CP-element group 57: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/$exit
      -- CP-element group 57: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/phi_stmt_1522/phi_stmt_1522_req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1522_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1522_req_4258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1522_req_4258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(57), ack => phi_stmt_1522_req_1); -- 
    sendB_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(55) & sendB_CP_3659_elements(56);
      gj_sendB_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	54 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1460/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    -- logger for CP element group sendB_CP_3659_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(58) fired."); 
        -- 
      end if; --
    end process; 
    sendB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(54) & sendB_CP_3659_elements(57);
      gj_sendB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	51 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_1460/merge_stmt_1514_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1460/merge_stmt_1514_PhiAck/$entry
      -- 
    -- logger for CP element group sendB_CP_3659_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(59) fired."); 
        -- 
      end if; --
    end process; 
    sendB_CP_3659_elements(59) <= OrReduce(sendB_CP_3659_elements(51) & sendB_CP_3659_elements(58));
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1460/merge_stmt_1514_PhiAck/phi_stmt_1515_ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1515_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1515_ack_4263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1515_ack_0, ack => sendB_CP_3659_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1460/merge_stmt_1514_PhiAck/phi_stmt_1522_ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1522_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1522_ack_4264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1522_ack_0, ack => sendB_CP_3659_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  place  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	8 
    -- CP-element group 62: 	9 
    -- CP-element group 62: 	11 
    -- CP-element group 62: 	13 
    -- CP-element group 62:  members (28) 
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/$entry
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_scale_1/scale_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_scale_1/scale_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_resized_1
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_scale_1/$entry
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_scale_1/$exit
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_scaled_1
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_computed_1
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_resize_1/$entry
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_resize_1/$exit
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_resize_1/index_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_index_resize_1/index_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1460/merge_stmt_1514__exit__
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556__entry__
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_final_index_sum_regn_update_start
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_final_index_sum_regn_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_final_index_sum_regn_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_final_index_sum_regn_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/array_obj_ref_1534_final_index_sum_regn_Update/req
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_complete/$entry
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/addr_of_1535_complete/req
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/word_access_complete/$entry
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/word_access_complete/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_1460/assign_stmt_1536_to_assign_stmt_1556/ptr_deref_1539_Update/word_access_complete/word_0/cr
      -- CP-element group 62: 	 branch_block_stmt_1460/merge_stmt_1514_PhiAck/$exit
      -- 
    -- logger for CP element group sendB_CP_3659_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:array_obj_ref_1534_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:array_obj_ref_1534_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:addr_of_1535_final_reg_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1539_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(62), ack => array_obj_ref_1534_index_offset_req_0); -- 
    req_3824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(62), ack => array_obj_ref_1534_index_offset_req_1); -- 
    req_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(62), ack => addr_of_1535_final_reg_req_1); -- 
    cr_3884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(62), ack => ptr_deref_1539_load_0_req_1); -- 
    sendB_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(60) & sendB_CP_3659_elements(61);
      gj_sendB_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	15 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/SplitProtocol/Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1567_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1567_inst_ack_0, ack => sendB_CP_3659_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	15 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/SplitProtocol/Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group sendB_CP_3659_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1567_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1567_inst_ack_1, ack => sendB_CP_3659_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	72 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/$exit
      -- CP-element group 65: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/$exit
      -- CP-element group 65: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/$exit
      -- CP-element group 65: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1567/SplitProtocol/$exit
      -- CP-element group 65: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1564/phi_stmt_1564_req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1564_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1564_req_4294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1564_req_4294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(65), ack => phi_stmt_1564_req_0); -- 
    sendB_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(63) & sendB_CP_3659_elements(64);
      gj_sendB_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	15 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/SplitProtocol/Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1571_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1571_inst_ack_0, ack => sendB_CP_3659_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	15 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/SplitProtocol/Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group sendB_CP_3659_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1571_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1571_inst_ack_1, ack => sendB_CP_3659_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	72 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/$exit
      -- CP-element group 68: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/$exit
      -- CP-element group 68: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/$exit
      -- CP-element group 68: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_sources/type_cast_1571/SplitProtocol/$exit
      -- CP-element group 68: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1568/phi_stmt_1568_req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1568_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1568_req_4317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1568_req_4317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(68), ack => phi_stmt_1568_req_0); -- 
    sendB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(66) & sendB_CP_3659_elements(67);
      gj_sendB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	15 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/SplitProtocol/Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1575_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1575_inst_ack_0, ack => sendB_CP_3659_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	15 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/SplitProtocol/Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group sendB_CP_3659_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1575_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1575_inst_ack_1, ack => sendB_CP_3659_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/$exit
      -- CP-element group 71: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/$exit
      -- CP-element group 71: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_sources/type_cast_1575/SplitProtocol/$exit
      -- CP-element group 71: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/phi_stmt_1572/phi_stmt_1572_req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1572_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1572_req_4340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1572_req_4340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(71), ack => phi_stmt_1572_req_0); -- 
    sendB_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(69) & sendB_CP_3659_elements(70);
      gj_sendB_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  join  fork  transition  place  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	65 
    -- CP-element group 72: 	68 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	74 
    -- CP-element group 72: 	75 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1460/forx_xbody_forx_xend_PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_1460/merge_stmt_1563_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1460/merge_stmt_1563_PhiAck/$entry
      -- 
    -- logger for CP element group sendB_CP_3659_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(72) fired."); 
        -- 
      end if; --
    end process; 
    sendB_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(65) & sendB_CP_3659_elements(68) & sendB_CP_3659_elements(71);
      gj_sendB_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	76 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1460/merge_stmt_1563_PhiAck/phi_stmt_1564_ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1564_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1564_ack_4345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1564_ack_0, ack => sendB_CP_3659_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1460/merge_stmt_1563_PhiAck/phi_stmt_1568_ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1568_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1568_ack_4346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1568_ack_0, ack => sendB_CP_3659_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	72 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1460/merge_stmt_1563_PhiAck/phi_stmt_1572_ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1572_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1572_ack_4347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1572_ack_0, ack => sendB_CP_3659_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	73 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	1 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1460/merge_stmt_1563_PhiAck/$exit
      -- 
    -- logger for CP element group sendB_CP_3659_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(76) fired."); 
        -- 
      end if; --
    end process; 
    sendB_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(73) & sendB_CP_3659_elements(74) & sendB_CP_3659_elements(75);
      gj_sendB_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	20 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_1460/bbx_xnph_forx_xbody15_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_1460/bbx_xnph_forx_xbody15_PhiReq/phi_stmt_1621/$exit
      -- CP-element group 77: 	 branch_block_stmt_1460/bbx_xnph_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_1460/bbx_xnph_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1625_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_1460/bbx_xnph_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1621_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1621_req_4370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1621_req_4370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(77), ack => phi_stmt_1621_req_0); -- 
    -- Element group sendB_CP_3659_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => sendB_CP_3659_elements(20), ack => sendB_CP_3659_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	48 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group sendB_CP_3659_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1627_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_0, ack => sendB_CP_3659_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	48 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group sendB_CP_3659_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1627_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_1, ack => sendB_CP_3659_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/$exit
      -- CP-element group 80: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/$exit
      -- CP-element group 80: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/$exit
      -- CP-element group 80: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_1460/forx_xbody15_forx_xbody15_PhiReq/phi_stmt_1621/phi_stmt_1621_req
      -- 
    -- logger for CP element group sendB_CP_3659_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1621_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1621_req_4396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1621_req_4396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(80), ack => phi_stmt_1621_req_1); -- 
    sendB_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_3659_elements(78) & sendB_CP_3659_elements(79);
      gj_sendB_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_3659_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  merge  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1460/merge_stmt_1620_PhiReqMerge
      -- CP-element group 81: 	 branch_block_stmt_1460/merge_stmt_1620_PhiAck/$entry
      -- 
    -- logger for CP element group sendB_CP_3659_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(81) fired."); 
        -- 
      end if; --
    end process; 
    sendB_CP_3659_elements(81) <= OrReduce(sendB_CP_3659_elements(77) & sendB_CP_3659_elements(80));
    -- CP-element group 82:  fork  transition  place  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	21 
    -- CP-element group 82: 	22 
    -- CP-element group 82: 	24 
    -- CP-element group 82: 	26 
    -- CP-element group 82: 	28 
    -- CP-element group 82: 	30 
    -- CP-element group 82: 	32 
    -- CP-element group 82: 	34 
    -- CP-element group 82:  members (41) 
      -- CP-element group 82: 	 branch_block_stmt_1460/merge_stmt_1620__exit__
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696__entry__
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_resized_1
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_scaled_1
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_computed_1
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_resize_1/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_resize_1/$exit
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_resize_1/index_resize_req
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_resize_1/index_resize_ack
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_scale_1/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_scale_1/$exit
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_scale_1/scale_rename_req
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_index_scale_1/scale_rename_ack
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_final_index_sum_regn_update_start
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_final_index_sum_regn_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_final_index_sum_regn_Sample/req
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_final_index_sum_regn_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/array_obj_ref_1633_final_index_sum_regn_Update/req
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_complete/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/addr_of_1634_complete/req
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/word_access_complete/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/word_access_complete/word_0/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/ptr_deref_1638_Update/word_access_complete/word_0/cr
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1642_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1652_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1662_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1460/assign_stmt_1635_to_assign_stmt_1696/type_cast_1672_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1460/merge_stmt_1620_PhiAck/$exit
      -- CP-element group 82: 	 branch_block_stmt_1460/merge_stmt_1620_PhiAck/phi_stmt_1621_ack
      -- 
    -- logger for CP element group sendB_CP_3659_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:phi_stmt_1621_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:array_obj_ref_1633_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:array_obj_ref_1633_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:addr_of_1634_final_reg_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:ptr_deref_1638_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1642_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1652_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1662_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:type_cast_1672_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1621_ack_4401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1621_ack_0, ack => sendB_CP_3659_elements(82)); -- 
    req_3976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(82), ack => array_obj_ref_1633_index_offset_req_0); -- 
    req_3981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(82), ack => array_obj_ref_1633_index_offset_req_1); -- 
    req_3996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(82), ack => addr_of_1634_final_reg_req_1); -- 
    cr_4041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(82), ack => ptr_deref_1638_load_0_req_1); -- 
    cr_4060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(82), ack => type_cast_1642_inst_req_1); -- 
    cr_4074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(82), ack => type_cast_1652_inst_req_1); -- 
    cr_4088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(82), ack => type_cast_1662_inst_req_1); -- 
    cr_4102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_3659_elements(82), ack => type_cast_1672_inst_req_1); -- 
    -- CP-element group 83:  merge  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	4 
    -- CP-element group 83: 	18 
    -- CP-element group 83: 	47 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (16) 
      -- CP-element group 83: 	 $exit
      -- CP-element group 83: 	 branch_block_stmt_1460/$exit
      -- CP-element group 83: 	 branch_block_stmt_1460/branch_block_stmt_1460__exit__
      -- CP-element group 83: 	 branch_block_stmt_1460/merge_stmt_1705__exit__
      -- CP-element group 83: 	 branch_block_stmt_1460/return__
      -- CP-element group 83: 	 branch_block_stmt_1460/merge_stmt_1707__exit__
      -- CP-element group 83: 	 branch_block_stmt_1460/merge_stmt_1705_PhiReqMerge
      -- CP-element group 83: 	 branch_block_stmt_1460/merge_stmt_1705_PhiAck/$entry
      -- CP-element group 83: 	 branch_block_stmt_1460/merge_stmt_1705_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_1460/merge_stmt_1705_PhiAck/dummy
      -- CP-element group 83: 	 branch_block_stmt_1460/return___PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_1460/return___PhiReq/$exit
      -- CP-element group 83: 	 branch_block_stmt_1460/merge_stmt_1707_PhiReqMerge
      -- CP-element group 83: 	 branch_block_stmt_1460/merge_stmt_1707_PhiAck/$entry
      -- CP-element group 83: 	 branch_block_stmt_1460/merge_stmt_1707_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_1460/merge_stmt_1707_PhiAck/dummy
      -- 
    -- logger for CP element group sendB_CP_3659_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and sendB_CP_3659_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:sendB:CP:sendB_CP_3659_elements(83) fired."); 
        -- 
      end if; --
    end process; 
    sendB_CP_3659_elements(83) <= OrReduce(sendB_CP_3659_elements(4) & sendB_CP_3659_elements(18) & sendB_CP_3659_elements(47));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar66_1533_resized : std_logic_vector(6 downto 0);
    signal R_indvar66_1533_scaled : std_logic_vector(6 downto 0);
    signal R_indvar_1632_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1632_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1534_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_1534_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_1534_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_1534_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_1534_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1534_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1633_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1633_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1633_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1633_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1633_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1633_root_address : std_logic_vector(13 downto 0);
    signal arrayidx19_1635 : std_logic_vector(31 downto 0);
    signal arrayidx_1536 : std_logic_vector(31 downto 0);
    signal cmp1357_1582 : std_logic_vector(0 downto 0);
    signal cmp60_1476 : std_logic_vector(0 downto 0);
    signal conv23_1643 : std_logic_vector(15 downto 0);
    signal conv29_1653 : std_logic_vector(15 downto 0);
    signal conv35_1663 : std_logic_vector(15 downto 0);
    signal conv41_1673 : std_logic_vector(15 downto 0);
    signal exitcond7_1696 : std_logic_vector(0 downto 0);
    signal exitcond_1556 : std_logic_vector(0 downto 0);
    signal iNsTr_0_1466 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1499 : std_logic_vector(63 downto 0);
    signal indvar66_1515 : std_logic_vector(63 downto 0);
    signal indvar_1621 : std_logic_vector(63 downto 0);
    signal indvarx_xnext67_1551 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1691 : std_logic_vector(63 downto 0);
    signal mul_1545 : std_logic_vector(31 downto 0);
    signal mulx_xlcssa_1564 : std_logic_vector(31 downto 0);
    signal num_elemsx_x061_1522 : std_logic_vector(31 downto 0);
    signal num_elemsx_x061x_xlcssa_1572 : std_logic_vector(31 downto 0);
    signal ptr_deref_1469_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1469_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1469_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1469_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1469_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1539_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1539_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1539_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1539_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1539_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1638_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1638_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1638_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1638_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1638_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr26_1649 : std_logic_vector(63 downto 0);
    signal shr32_1659 : std_logic_vector(63 downto 0);
    signal shr38_1669 : std_logic_vector(63 downto 0);
    signal tmp159_1470 : std_logic_vector(31 downto 0);
    signal tmp1_1594 : std_logic_vector(31 downto 0);
    signal tmp1x_xop_1495 : std_logic_vector(31 downto 0);
    signal tmp20_1639 : std_logic_vector(63 downto 0);
    signal tmp2_1599 : std_logic_vector(63 downto 0);
    signal tmp3_1540 : std_logic_vector(31 downto 0);
    signal tmp3x_xlcssa_1568 : std_logic_vector(31 downto 0);
    signal tmp4_1605 : std_logic_vector(63 downto 0);
    signal tmp5_1611 : std_logic_vector(0 downto 0);
    signal tmp68_1489 : std_logic_vector(0 downto 0);
    signal tmp72_1512 : std_logic_vector(63 downto 0);
    signal type_cast_1474_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1487_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1493_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1503_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1510_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1519_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1521_wire : std_logic_vector(63 downto 0);
    signal type_cast_1526_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1528_wire : std_logic_vector(31 downto 0);
    signal type_cast_1549_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1567_wire : std_logic_vector(31 downto 0);
    signal type_cast_1571_wire : std_logic_vector(31 downto 0);
    signal type_cast_1575_wire : std_logic_vector(31 downto 0);
    signal type_cast_1580_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1597_wire : std_logic_vector(63 downto 0);
    signal type_cast_1603_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1609_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1616_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1625_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1627_wire : std_logic_vector(63 downto 0);
    signal type_cast_1647_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1657_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1667_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1689_wire_constant : std_logic_vector(63 downto 0);
    signal umax6_1618 : std_logic_vector(63 downto 0);
    signal xx_xop_1505 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1534_constant_part_of_offset <= "0000010";
    array_obj_ref_1534_offset_scale_factor_0 <= "1000000";
    array_obj_ref_1534_offset_scale_factor_1 <= "0000001";
    array_obj_ref_1534_resized_base_address <= "0000000";
    array_obj_ref_1633_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1633_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1633_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1633_resized_base_address <= "00000000000000";
    iNsTr_0_1466 <= "00000000000000000000000000000001";
    ptr_deref_1469_word_offset_0 <= "0000000";
    ptr_deref_1539_word_offset_0 <= "0000000";
    ptr_deref_1638_word_offset_0 <= "00000000000000";
    type_cast_1474_wire_constant <= "00000000000000000000000000000000";
    type_cast_1487_wire_constant <= "00000000000000000000000000000001";
    type_cast_1493_wire_constant <= "11111111111111111111111111111111";
    type_cast_1503_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1510_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1519_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1526_wire_constant <= "00000000000000000000000000000001";
    type_cast_1549_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1580_wire_constant <= "00000000000000000000000000000011";
    type_cast_1603_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1609_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1616_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1625_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1647_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1657_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1667_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1689_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    -- logger for phi phi_stmt_1515
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1515_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:sendB:DP:phi_stmt_1515:input-0 type_cast_1519_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1519_wire_constant));
          --
        end if;
        if phi_stmt_1515_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:sendB:DP:phi_stmt_1515:input-1 type_cast_1521_wire= " & Convert_SLV_To_Hex_String(type_cast_1521_wire));
          --
        end if;
        if phi_stmt_1515_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:sendB:DP:phi_stmt_1515:sample-completed");
          --
        end if;
        if phi_stmt_1515_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:sendB:DP:phi_stmt_1515:output indvar66_1515= " & Convert_SLV_To_Hex_String(indvar66_1515));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1515: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1519_wire_constant & type_cast_1521_wire;
      req <= phi_stmt_1515_req_0 & phi_stmt_1515_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1515",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1515_ack_0,
          idata => idata,
          odata => indvar66_1515,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1515
    -- logger for phi phi_stmt_1522
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1522_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:sendB:DP:phi_stmt_1522:input-0 type_cast_1526_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1526_wire_constant));
          --
        end if;
        if phi_stmt_1522_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:sendB:DP:phi_stmt_1522:input-1 type_cast_1528_wire= " & Convert_SLV_To_Hex_String(type_cast_1528_wire));
          --
        end if;
        if phi_stmt_1522_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:sendB:DP:phi_stmt_1522:sample-completed");
          --
        end if;
        if phi_stmt_1522_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:sendB:DP:phi_stmt_1522:output num_elemsx_x061_1522= " & Convert_SLV_To_Hex_String(num_elemsx_x061_1522));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1522: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1526_wire_constant & type_cast_1528_wire;
      req <= phi_stmt_1522_req_0 & phi_stmt_1522_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1522",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1522_ack_0,
          idata => idata,
          odata => num_elemsx_x061_1522,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1522
    -- logger for phi phi_stmt_1564
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1564_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:sendB:DP:phi_stmt_1564:input-0 type_cast_1567_wire= " & Convert_SLV_To_Hex_String(type_cast_1567_wire));
          --
        end if;
        if phi_stmt_1564_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:sendB:DP:phi_stmt_1564:sample-completed");
          --
        end if;
        if phi_stmt_1564_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:sendB:DP:phi_stmt_1564:output mulx_xlcssa_1564= " & Convert_SLV_To_Hex_String(mulx_xlcssa_1564));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1564: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1567_wire;
      req(0) <= phi_stmt_1564_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1564",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1564_ack_0,
          idata => idata,
          odata => mulx_xlcssa_1564,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1564
    -- logger for phi phi_stmt_1568
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1568_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:sendB:DP:phi_stmt_1568:input-0 type_cast_1571_wire= " & Convert_SLV_To_Hex_String(type_cast_1571_wire));
          --
        end if;
        if phi_stmt_1568_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:sendB:DP:phi_stmt_1568:sample-completed");
          --
        end if;
        if phi_stmt_1568_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:sendB:DP:phi_stmt_1568:output tmp3x_xlcssa_1568= " & Convert_SLV_To_Hex_String(tmp3x_xlcssa_1568));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1568: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1571_wire;
      req(0) <= phi_stmt_1568_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1568",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1568_ack_0,
          idata => idata,
          odata => tmp3x_xlcssa_1568,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1568
    -- logger for phi phi_stmt_1572
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1572_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:sendB:DP:phi_stmt_1572:input-0 type_cast_1575_wire= " & Convert_SLV_To_Hex_String(type_cast_1575_wire));
          --
        end if;
        if phi_stmt_1572_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:sendB:DP:phi_stmt_1572:sample-completed");
          --
        end if;
        if phi_stmt_1572_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:sendB:DP:phi_stmt_1572:output num_elemsx_x061x_xlcssa_1572= " & Convert_SLV_To_Hex_String(num_elemsx_x061x_xlcssa_1572));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1572: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1575_wire;
      req(0) <= phi_stmt_1572_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1572",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1572_ack_0,
          idata => idata,
          odata => num_elemsx_x061x_xlcssa_1572,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1572
    -- logger for phi phi_stmt_1621
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1621_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:sendB:DP:phi_stmt_1621:input-0 type_cast_1625_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1625_wire_constant));
          --
        end if;
        if phi_stmt_1621_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:sendB:DP:phi_stmt_1621:input-1 type_cast_1627_wire= " & Convert_SLV_To_Hex_String(type_cast_1627_wire));
          --
        end if;
        if phi_stmt_1621_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:sendB:DP:phi_stmt_1621:sample-completed");
          --
        end if;
        if phi_stmt_1621_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:sendB:DP:phi_stmt_1621:output indvar_1621= " & Convert_SLV_To_Hex_String(indvar_1621));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1621: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1625_wire_constant & type_cast_1627_wire;
      req <= phi_stmt_1621_req_0 & phi_stmt_1621_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1621",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1621_ack_0,
          idata => idata,
          odata => indvar_1621,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1621
    -- logger for split-operator MUX_1511_inst flow-through 
    process(tmp72_1512) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:MUX_1511_inst:flowthrough inputs: " & " tmp68_1489 = "& Convert_SLV_To_Hex_String(tmp68_1489) & " xx_xop_1505 = "& Convert_SLV_To_Hex_String(xx_xop_1505) & " type_cast_1510_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1510_wire_constant) & " outputs:" & " tmp72_1512= "  & Convert_SLV_To_Hex_String(tmp72_1512));
      --
    end process; 
    -- flow-through select operator MUX_1511_inst
    tmp72_1512 <= xx_xop_1505 when (tmp68_1489(0) /=  '0') else type_cast_1510_wire_constant;
    -- logger for split-operator MUX_1617_inst flow-through 
    process(umax6_1618) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:MUX_1617_inst:flowthrough inputs: " & " tmp5_1611 = "& Convert_SLV_To_Hex_String(tmp5_1611) & " tmp4_1605 = "& Convert_SLV_To_Hex_String(tmp4_1605) & " type_cast_1616_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1616_wire_constant) & " outputs:" & " umax6_1618= "  & Convert_SLV_To_Hex_String(umax6_1618));
      --
    end process; 
    -- flow-through select operator MUX_1617_inst
    umax6_1618 <= tmp4_1605 when (tmp5_1611(0) /=  '0') else type_cast_1616_wire_constant;
    -- logger for split-operator addr_of_1535_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_1535_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:addr_of_1535_final_reg:started:   inputs: " & " array_obj_ref_1534_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1534_root_address));
          --
        end if; 
        if addr_of_1535_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:addr_of_1535_final_reg:finished:  outputs: " & " arrayidx_1536= "  & Convert_SLV_To_Hex_String(arrayidx_1536));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_1535_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1535_final_reg_req_0;
      addr_of_1535_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1535_final_reg_req_1;
      addr_of_1535_final_reg_ack_1<= rack(0);
      addr_of_1535_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1535_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1534_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1536,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_1634_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_1634_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:addr_of_1634_final_reg:started:   inputs: " & " array_obj_ref_1633_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1633_root_address));
          --
        end if; 
        if addr_of_1634_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:addr_of_1634_final_reg:finished:  outputs: " & " arrayidx19_1635= "  & Convert_SLV_To_Hex_String(arrayidx19_1635));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_1634_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1634_final_reg_req_0;
      addr_of_1634_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1634_final_reg_req_1;
      addr_of_1634_final_reg_ack_1<= rack(0);
      addr_of_1634_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1634_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1633_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx19_1635,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1498_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1498_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1498_inst:started:   inputs: " & " tmp1x_xop_1495 = "& Convert_SLV_To_Hex_String(tmp1x_xop_1495));
          --
        end if; 
        if type_cast_1498_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1498_inst:finished:  outputs: " & " iNsTr_3_1499= "  & Convert_SLV_To_Hex_String(iNsTr_3_1499));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1498_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1498_inst_req_0;
      type_cast_1498_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1498_inst_req_1;
      type_cast_1498_inst_ack_1<= rack(0);
      type_cast_1498_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1498_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1x_xop_1495,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_3_1499,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1521_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1521_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1521_inst:started:   inputs: " & " indvarx_xnext67_1551 = "& Convert_SLV_To_Hex_String(indvarx_xnext67_1551));
          --
        end if; 
        if type_cast_1521_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1521_inst:finished:  outputs: " & " type_cast_1521_wire= "  & Convert_SLV_To_Hex_String(type_cast_1521_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1521_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1521_inst_req_0;
      type_cast_1521_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1521_inst_req_1;
      type_cast_1521_inst_ack_1<= rack(0);
      type_cast_1521_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1521_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext67_1551,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1521_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1528_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1528_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1528_inst:started:   inputs: " & " mul_1545 = "& Convert_SLV_To_Hex_String(mul_1545));
          --
        end if; 
        if type_cast_1528_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1528_inst:finished:  outputs: " & " type_cast_1528_wire= "  & Convert_SLV_To_Hex_String(type_cast_1528_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1528_inst_req_0;
      type_cast_1528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1528_inst_req_1;
      type_cast_1528_inst_ack_1<= rack(0);
      type_cast_1528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul_1545,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1528_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1567_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1567_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1567_inst:started:   inputs: " & " mul_1545 = "& Convert_SLV_To_Hex_String(mul_1545));
          --
        end if; 
        if type_cast_1567_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1567_inst:finished:  outputs: " & " type_cast_1567_wire= "  & Convert_SLV_To_Hex_String(type_cast_1567_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1567_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1567_inst_req_0;
      type_cast_1567_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1567_inst_req_1;
      type_cast_1567_inst_ack_1<= rack(0);
      type_cast_1567_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1567_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul_1545,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1567_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1571_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1571_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1571_inst:started:   inputs: " & " tmp3_1540 = "& Convert_SLV_To_Hex_String(tmp3_1540));
          --
        end if; 
        if type_cast_1571_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1571_inst:finished:  outputs: " & " type_cast_1571_wire= "  & Convert_SLV_To_Hex_String(type_cast_1571_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1571_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1571_inst_req_0;
      type_cast_1571_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1571_inst_req_1;
      type_cast_1571_inst_ack_1<= rack(0);
      type_cast_1571_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1571_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_1540,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1571_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1575_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1575_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1575_inst:started:   inputs: " & " num_elemsx_x061_1522 = "& Convert_SLV_To_Hex_String(num_elemsx_x061_1522));
          --
        end if; 
        if type_cast_1575_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1575_inst:finished:  outputs: " & " type_cast_1575_wire= "  & Convert_SLV_To_Hex_String(type_cast_1575_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1575_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1575_inst_req_0;
      type_cast_1575_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1575_inst_req_1;
      type_cast_1575_inst_ack_1<= rack(0);
      type_cast_1575_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1575_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_elemsx_x061_1522,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1575_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1598_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1598_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1598_inst:started:   inputs: " & " type_cast_1597_wire = "& Convert_SLV_To_Hex_String(type_cast_1597_wire));
          --
        end if; 
        if type_cast_1598_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1598_inst:finished:  outputs: " & " tmp2_1599= "  & Convert_SLV_To_Hex_String(tmp2_1599));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1598_inst_req_0;
      type_cast_1598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1598_inst_req_1;
      type_cast_1598_inst_ack_1<= rack(0);
      type_cast_1598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1597_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp2_1599,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1627_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1627_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1627_inst:started:   inputs: " & " indvarx_xnext_1691 = "& Convert_SLV_To_Hex_String(indvarx_xnext_1691));
          --
        end if; 
        if type_cast_1627_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1627_inst:finished:  outputs: " & " type_cast_1627_wire= "  & Convert_SLV_To_Hex_String(type_cast_1627_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1627_inst_req_0;
      type_cast_1627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1627_inst_req_1;
      type_cast_1627_inst_ack_1<= rack(0);
      type_cast_1627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1691,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1627_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1642_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1642_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1642_inst:started:   inputs: " & " tmp20_1639 = "& Convert_SLV_To_Hex_String(tmp20_1639));
          --
        end if; 
        if type_cast_1642_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1642_inst:finished:  outputs: " & " conv23_1643= "  & Convert_SLV_To_Hex_String(conv23_1643));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1642_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1642_inst_req_0;
      type_cast_1642_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1642_inst_req_1;
      type_cast_1642_inst_ack_1<= rack(0);
      type_cast_1642_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1642_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp20_1639,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_1643,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1652_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1652_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1652_inst:started:   inputs: " & " shr26_1649 = "& Convert_SLV_To_Hex_String(shr26_1649));
          --
        end if; 
        if type_cast_1652_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1652_inst:finished:  outputs: " & " conv29_1653= "  & Convert_SLV_To_Hex_String(conv29_1653));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1652_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1652_inst_req_0;
      type_cast_1652_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1652_inst_req_1;
      type_cast_1652_inst_ack_1<= rack(0);
      type_cast_1652_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1652_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr26_1649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1653,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1662_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1662_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1662_inst:started:   inputs: " & " shr32_1659 = "& Convert_SLV_To_Hex_String(shr32_1659));
          --
        end if; 
        if type_cast_1662_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1662_inst:finished:  outputs: " & " conv35_1663= "  & Convert_SLV_To_Hex_String(conv35_1663));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1662_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1662_inst_req_0;
      type_cast_1662_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1662_inst_req_1;
      type_cast_1662_inst_ack_1<= rack(0);
      type_cast_1662_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1662_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr32_1659,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_1663,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1672_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1672_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1672_inst:started:   inputs: " & " shr38_1669 = "& Convert_SLV_To_Hex_String(shr38_1669));
          --
        end if; 
        if type_cast_1672_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1672_inst:finished:  outputs: " & " conv41_1673= "  & Convert_SLV_To_Hex_String(conv41_1673));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1672_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1672_inst_req_0;
      type_cast_1672_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1672_inst_req_1;
      type_cast_1672_inst_ack_1<= rack(0);
      type_cast_1672_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1672_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr38_1669,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_1673,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_1534_index_1_rename flow-through 
    process(R_indvar66_1533_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:array_obj_ref_1534_index_1_rename:flowthrough  inputs: " & " R_indvar66_1533_resized = "& Convert_SLV_To_Hex_String(R_indvar66_1533_resized) & "outputs: " & " R_indvar66_1533_scaled= "  & Convert_SLV_To_Hex_String(R_indvar66_1533_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1534_index_1_rename
    process(R_indvar66_1533_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar66_1533_resized;
      ov(6 downto 0) := iv;
      R_indvar66_1533_scaled <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1534_index_1_resize flow-through 
    process(R_indvar66_1533_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:array_obj_ref_1534_index_1_resize:flowthrough  inputs: " & " indvar66_1515 = "& Convert_SLV_To_Hex_String(indvar66_1515) & "outputs: " & " R_indvar66_1533_resized= "  & Convert_SLV_To_Hex_String(R_indvar66_1533_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1534_index_1_resize
    process(indvar66_1515) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar66_1515;
      ov := iv(6 downto 0);
      R_indvar66_1533_resized <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1534_root_address_inst flow-through 
    process(array_obj_ref_1534_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:array_obj_ref_1534_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1534_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1534_final_offset) & "outputs: " & " array_obj_ref_1534_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1534_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1534_root_address_inst
    process(array_obj_ref_1534_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1534_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_1534_root_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1633_index_1_rename flow-through 
    process(R_indvar_1632_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:array_obj_ref_1633_index_1_rename:flowthrough  inputs: " & " R_indvar_1632_resized = "& Convert_SLV_To_Hex_String(R_indvar_1632_resized) & "outputs: " & " R_indvar_1632_scaled= "  & Convert_SLV_To_Hex_String(R_indvar_1632_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1633_index_1_rename
    process(R_indvar_1632_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1632_resized;
      ov(13 downto 0) := iv;
      R_indvar_1632_scaled <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1633_index_1_resize flow-through 
    process(R_indvar_1632_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:array_obj_ref_1633_index_1_resize:flowthrough  inputs: " & " indvar_1621 = "& Convert_SLV_To_Hex_String(indvar_1621) & "outputs: " & " R_indvar_1632_resized= "  & Convert_SLV_To_Hex_String(R_indvar_1632_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1633_index_1_resize
    process(indvar_1621) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1621;
      ov := iv(13 downto 0);
      R_indvar_1632_resized <= ov(13 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1633_root_address_inst flow-through 
    process(array_obj_ref_1633_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:array_obj_ref_1633_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1633_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1633_final_offset) & "outputs: " & " array_obj_ref_1633_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1633_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1633_root_address_inst
    process(array_obj_ref_1633_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1633_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1633_root_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1469_addr_0 flow-through 
    process(ptr_deref_1469_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1469_addr_0:flowthrough  inputs: " & " ptr_deref_1469_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1469_root_address) & "outputs: " & " ptr_deref_1469_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1469_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1469_addr_0
    process(ptr_deref_1469_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1469_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1469_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1469_base_resize flow-through 
    process(ptr_deref_1469_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1469_base_resize:flowthrough  inputs: " & " iNsTr_0_1466 = "& Convert_SLV_To_Hex_String(iNsTr_0_1466) & "outputs: " & " ptr_deref_1469_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1469_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1469_base_resize
    process(iNsTr_0_1466) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_1466;
      ov := iv(6 downto 0);
      ptr_deref_1469_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1469_gather_scatter flow-through 
    process(tmp159_1470) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1469_gather_scatter:flowthrough  inputs: " & " ptr_deref_1469_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1469_data_0) & "outputs: " & " tmp159_1470= "  & Convert_SLV_To_Hex_String(tmp159_1470));
      --
    end process; 
    -- equivalence ptr_deref_1469_gather_scatter
    process(ptr_deref_1469_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1469_data_0;
      ov(31 downto 0) := iv;
      tmp159_1470 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1469_root_address_inst flow-through 
    process(ptr_deref_1469_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1469_root_address_inst:flowthrough  inputs: " & " ptr_deref_1469_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1469_resized_base_address) & "outputs: " & " ptr_deref_1469_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1469_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1469_root_address_inst
    process(ptr_deref_1469_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1469_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1469_root_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1539_addr_0 flow-through 
    process(ptr_deref_1539_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1539_addr_0:flowthrough  inputs: " & " ptr_deref_1539_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1539_root_address) & "outputs: " & " ptr_deref_1539_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1539_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1539_addr_0
    process(ptr_deref_1539_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1539_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1539_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1539_base_resize flow-through 
    process(ptr_deref_1539_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1539_base_resize:flowthrough  inputs: " & " arrayidx_1536 = "& Convert_SLV_To_Hex_String(arrayidx_1536) & "outputs: " & " ptr_deref_1539_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1539_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1539_base_resize
    process(arrayidx_1536) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1536;
      ov := iv(6 downto 0);
      ptr_deref_1539_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1539_gather_scatter flow-through 
    process(tmp3_1540) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1539_gather_scatter:flowthrough  inputs: " & " ptr_deref_1539_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1539_data_0) & "outputs: " & " tmp3_1540= "  & Convert_SLV_To_Hex_String(tmp3_1540));
      --
    end process; 
    -- equivalence ptr_deref_1539_gather_scatter
    process(ptr_deref_1539_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1539_data_0;
      ov(31 downto 0) := iv;
      tmp3_1540 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1539_root_address_inst flow-through 
    process(ptr_deref_1539_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1539_root_address_inst:flowthrough  inputs: " & " ptr_deref_1539_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1539_resized_base_address) & "outputs: " & " ptr_deref_1539_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1539_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1539_root_address_inst
    process(ptr_deref_1539_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1539_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1539_root_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1638_addr_0 flow-through 
    process(ptr_deref_1638_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1638_addr_0:flowthrough  inputs: " & " ptr_deref_1638_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_1638_root_address) & "outputs: " & " ptr_deref_1638_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1638_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_1638_addr_0
    process(ptr_deref_1638_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1638_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1638_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1638_base_resize flow-through 
    process(ptr_deref_1638_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1638_base_resize:flowthrough  inputs: " & " arrayidx19_1635 = "& Convert_SLV_To_Hex_String(arrayidx19_1635) & "outputs: " & " ptr_deref_1638_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1638_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_1638_base_resize
    process(arrayidx19_1635) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx19_1635;
      ov := iv(13 downto 0);
      ptr_deref_1638_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1638_gather_scatter flow-through 
    process(tmp20_1639) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1638_gather_scatter:flowthrough  inputs: " & " ptr_deref_1638_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1638_data_0) & "outputs: " & " tmp20_1639= "  & Convert_SLV_To_Hex_String(tmp20_1639));
      --
    end process; 
    -- equivalence ptr_deref_1638_gather_scatter
    process(ptr_deref_1638_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1638_data_0;
      ov(63 downto 0) := iv;
      tmp20_1639 <= ov(63 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_1638_root_address_inst flow-through 
    process(ptr_deref_1638_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1638_root_address_inst:flowthrough  inputs: " & " ptr_deref_1638_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_1638_resized_base_address) & "outputs: " & " ptr_deref_1638_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_1638_root_address));
      --
    end process; 
    -- equivalence ptr_deref_1638_root_address_inst
    process(ptr_deref_1638_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1638_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1638_root_address <= ov(13 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1477_branch_req_0," req0 if_stmt_1477_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1477_branch_ack_0," ack0 if_stmt_1477_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1477_branch_ack_1," ack1 if_stmt_1477_branch");
    if_stmt_1477_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp60_1476;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1477_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1477_branch_req_0,
          ack0 => if_stmt_1477_branch_ack_0,
          ack1 => if_stmt_1477_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1557_branch_req_0," req0 if_stmt_1557_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1557_branch_ack_0," ack0 if_stmt_1557_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1557_branch_ack_1," ack1 if_stmt_1557_branch");
    if_stmt_1557_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1556;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1557_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1557_branch_req_0,
          ack0 => if_stmt_1557_branch_ack_0,
          ack1 => if_stmt_1557_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1583_branch_req_0," req0 if_stmt_1583_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1583_branch_ack_0," ack0 if_stmt_1583_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1583_branch_ack_1," ack1 if_stmt_1583_branch");
    if_stmt_1583_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1357_1582;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1583_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1583_branch_req_0,
          ack0 => if_stmt_1583_branch_ack_0,
          ack1 => if_stmt_1583_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1697_branch_req_0," req0 if_stmt_1697_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1697_branch_ack_0," ack0 if_stmt_1697_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1697_branch_ack_1," ack1 if_stmt_1697_branch");
    if_stmt_1697_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond7_1696;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1697_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1697_branch_req_0,
          ack0 => if_stmt_1697_branch_ack_0,
          ack1 => if_stmt_1697_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u32_u32_1494_inst flow-through 
    process(tmp1x_xop_1495) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ADD_u32_u32_1494_inst:flowthrough inputs: " & " tmp159_1470 = "& Convert_SLV_To_Hex_String(tmp159_1470) & " type_cast_1493_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1493_wire_constant) & " outputs:" & " tmp1x_xop_1495= "  & Convert_SLV_To_Hex_String(tmp1x_xop_1495));
      --
    end process; 
    -- binary operator ADD_u32_u32_1494_inst
    process(tmp159_1470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp159_1470, type_cast_1493_wire_constant, tmp_var);
      tmp1x_xop_1495 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_1504_inst flow-through 
    process(xx_xop_1505) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ADD_u64_u64_1504_inst:flowthrough inputs: " & " iNsTr_3_1499 = "& Convert_SLV_To_Hex_String(iNsTr_3_1499) & " type_cast_1503_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1503_wire_constant) & " outputs:" & " xx_xop_1505= "  & Convert_SLV_To_Hex_String(xx_xop_1505));
      --
    end process; 
    -- binary operator ADD_u64_u64_1504_inst
    process(iNsTr_3_1499) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_3_1499, type_cast_1503_wire_constant, tmp_var);
      xx_xop_1505 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_1550_inst flow-through 
    process(indvarx_xnext67_1551) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ADD_u64_u64_1550_inst:flowthrough inputs: " & " indvar66_1515 = "& Convert_SLV_To_Hex_String(indvar66_1515) & " type_cast_1549_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1549_wire_constant) & " outputs:" & " indvarx_xnext67_1551= "  & Convert_SLV_To_Hex_String(indvarx_xnext67_1551));
      --
    end process; 
    -- binary operator ADD_u64_u64_1550_inst
    process(indvar66_1515) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar66_1515, type_cast_1549_wire_constant, tmp_var);
      indvarx_xnext67_1551 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_1690_inst flow-through 
    process(indvarx_xnext_1691) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ADD_u64_u64_1690_inst:flowthrough inputs: " & " indvar_1621 = "& Convert_SLV_To_Hex_String(indvar_1621) & " type_cast_1689_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1689_wire_constant) & " outputs:" & " indvarx_xnext_1691= "  & Convert_SLV_To_Hex_String(indvarx_xnext_1691));
      --
    end process; 
    -- binary operator ADD_u64_u64_1690_inst
    process(indvar_1621) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1621, type_cast_1689_wire_constant, tmp_var);
      indvarx_xnext_1691 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u32_u1_1475_inst flow-through 
    process(cmp60_1476) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:EQ_u32_u1_1475_inst:flowthrough inputs: " & " tmp159_1470 = "& Convert_SLV_To_Hex_String(tmp159_1470) & " type_cast_1474_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1474_wire_constant) & " outputs:" & " cmp60_1476= "  & Convert_SLV_To_Hex_String(cmp60_1476));
      --
    end process; 
    -- binary operator EQ_u32_u1_1475_inst
    process(tmp159_1470) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tmp159_1470, type_cast_1474_wire_constant, tmp_var);
      cmp60_1476 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_1555_inst flow-through 
    process(exitcond_1556) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:EQ_u64_u1_1555_inst:flowthrough inputs: " & " indvarx_xnext67_1551 = "& Convert_SLV_To_Hex_String(indvarx_xnext67_1551) & " tmp72_1512 = "& Convert_SLV_To_Hex_String(tmp72_1512) & " outputs:" & " exitcond_1556= "  & Convert_SLV_To_Hex_String(exitcond_1556));
      --
    end process; 
    -- binary operator EQ_u64_u1_1555_inst
    process(indvarx_xnext67_1551, tmp72_1512) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext67_1551, tmp72_1512, tmp_var);
      exitcond_1556 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_1695_inst flow-through 
    process(exitcond7_1696) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:EQ_u64_u1_1695_inst:flowthrough inputs: " & " indvarx_xnext_1691 = "& Convert_SLV_To_Hex_String(indvarx_xnext_1691) & " umax6_1618 = "& Convert_SLV_To_Hex_String(umax6_1618) & " outputs:" & " exitcond7_1696= "  & Convert_SLV_To_Hex_String(exitcond7_1696));
      --
    end process; 
    -- binary operator EQ_u64_u1_1695_inst
    process(indvarx_xnext_1691, umax6_1618) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1691, umax6_1618, tmp_var);
      exitcond7_1696 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_1604_inst flow-through 
    process(tmp4_1605) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:LSHR_u64_u64_1604_inst:flowthrough inputs: " & " tmp2_1599 = "& Convert_SLV_To_Hex_String(tmp2_1599) & " type_cast_1603_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1603_wire_constant) & " outputs:" & " tmp4_1605= "  & Convert_SLV_To_Hex_String(tmp4_1605));
      --
    end process; 
    -- binary operator LSHR_u64_u64_1604_inst
    process(tmp2_1599) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_1599, type_cast_1603_wire_constant, tmp_var);
      tmp4_1605 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_1648_inst flow-through 
    process(shr26_1649) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:LSHR_u64_u64_1648_inst:flowthrough inputs: " & " tmp20_1639 = "& Convert_SLV_To_Hex_String(tmp20_1639) & " type_cast_1647_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1647_wire_constant) & " outputs:" & " shr26_1649= "  & Convert_SLV_To_Hex_String(shr26_1649));
      --
    end process; 
    -- binary operator LSHR_u64_u64_1648_inst
    process(tmp20_1639) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp20_1639, type_cast_1647_wire_constant, tmp_var);
      shr26_1649 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_1658_inst flow-through 
    process(shr32_1659) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:LSHR_u64_u64_1658_inst:flowthrough inputs: " & " tmp20_1639 = "& Convert_SLV_To_Hex_String(tmp20_1639) & " type_cast_1657_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1657_wire_constant) & " outputs:" & " shr32_1659= "  & Convert_SLV_To_Hex_String(shr32_1659));
      --
    end process; 
    -- binary operator LSHR_u64_u64_1658_inst
    process(tmp20_1639) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp20_1639, type_cast_1657_wire_constant, tmp_var);
      shr32_1659 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_1668_inst flow-through 
    process(shr38_1669) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:LSHR_u64_u64_1668_inst:flowthrough inputs: " & " tmp20_1639 = "& Convert_SLV_To_Hex_String(tmp20_1639) & " type_cast_1667_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1667_wire_constant) & " outputs:" & " shr38_1669= "  & Convert_SLV_To_Hex_String(shr38_1669));
      --
    end process; 
    -- binary operator LSHR_u64_u64_1668_inst
    process(tmp20_1639) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp20_1639, type_cast_1667_wire_constant, tmp_var);
      shr38_1669 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_1544_inst flow-through 
    process(mul_1545) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:MUL_u32_u32_1544_inst:flowthrough inputs: " & " tmp3_1540 = "& Convert_SLV_To_Hex_String(tmp3_1540) & " num_elemsx_x061_1522 = "& Convert_SLV_To_Hex_String(num_elemsx_x061_1522) & " outputs:" & " mul_1545= "  & Convert_SLV_To_Hex_String(mul_1545));
      --
    end process; 
    -- binary operator MUL_u32_u32_1544_inst
    process(tmp3_1540, num_elemsx_x061_1522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp3_1540, num_elemsx_x061_1522, tmp_var);
      mul_1545 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_1593_inst flow-through 
    process(tmp1_1594) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:MUL_u32_u32_1593_inst:flowthrough inputs: " & " num_elemsx_x061x_xlcssa_1572 = "& Convert_SLV_To_Hex_String(num_elemsx_x061x_xlcssa_1572) & " tmp3x_xlcssa_1568 = "& Convert_SLV_To_Hex_String(tmp3x_xlcssa_1568) & " outputs:" & " tmp1_1594= "  & Convert_SLV_To_Hex_String(tmp1_1594));
      --
    end process; 
    -- binary operator MUL_u32_u32_1593_inst
    process(num_elemsx_x061x_xlcssa_1572, tmp3x_xlcssa_1568) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(num_elemsx_x061x_xlcssa_1572, tmp3x_xlcssa_1568, tmp_var);
      tmp1_1594 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u32_u1_1488_inst flow-through 
    process(tmp68_1489) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:UGT_u32_u1_1488_inst:flowthrough inputs: " & " tmp159_1470 = "& Convert_SLV_To_Hex_String(tmp159_1470) & " type_cast_1487_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1487_wire_constant) & " outputs:" & " tmp68_1489= "  & Convert_SLV_To_Hex_String(tmp68_1489));
      --
    end process; 
    -- binary operator UGT_u32_u1_1488_inst
    process(tmp159_1470) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp159_1470, type_cast_1487_wire_constant, tmp_var);
      tmp68_1489 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u32_u1_1581_inst flow-through 
    process(cmp1357_1582) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:UGT_u32_u1_1581_inst:flowthrough inputs: " & " mulx_xlcssa_1564 = "& Convert_SLV_To_Hex_String(mulx_xlcssa_1564) & " type_cast_1580_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1580_wire_constant) & " outputs:" & " cmp1357_1582= "  & Convert_SLV_To_Hex_String(cmp1357_1582));
      --
    end process; 
    -- binary operator UGT_u32_u1_1581_inst
    process(mulx_xlcssa_1564) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mulx_xlcssa_1564, type_cast_1580_wire_constant, tmp_var);
      cmp1357_1582 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u64_u1_1610_inst flow-through 
    process(tmp5_1611) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:UGT_u64_u1_1610_inst:flowthrough inputs: " & " tmp4_1605 = "& Convert_SLV_To_Hex_String(tmp4_1605) & " type_cast_1609_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1609_wire_constant) & " outputs:" & " tmp5_1611= "  & Convert_SLV_To_Hex_String(tmp5_1611));
      --
    end process; 
    -- binary operator UGT_u64_u1_1610_inst
    process(tmp4_1605) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp4_1605, type_cast_1609_wire_constant, tmp_var);
      tmp5_1611 <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_1534_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1534_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:array_obj_ref_1534_index_offset:started:   inputs: " & " R_indvar66_1533_scaled = "& Convert_SLV_To_Hex_String(R_indvar66_1533_scaled) & " array_obj_ref_1534_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1534_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1534_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:array_obj_ref_1534_index_offset:finished:  outputs: " & " array_obj_ref_1534_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1534_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (16) : array_obj_ref_1534_index_offset 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar66_1533_scaled;
      array_obj_ref_1534_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1534_index_offset_req_0;
      array_obj_ref_1534_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1534_index_offset_req_1;
      array_obj_ref_1534_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000010",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- logger for split-operator array_obj_ref_1633_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1633_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:array_obj_ref_1633_index_offset:started:   inputs: " & " R_indvar_1632_scaled = "& Convert_SLV_To_Hex_String(R_indvar_1632_scaled) & " array_obj_ref_1633_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1633_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1633_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:array_obj_ref_1633_index_offset:finished:  outputs: " & " array_obj_ref_1633_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1633_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (17) : array_obj_ref_1633_index_offset 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1632_scaled;
      array_obj_ref_1633_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1633_index_offset_req_0;
      array_obj_ref_1633_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1633_index_offset_req_1;
      array_obj_ref_1633_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- logger for split-operator type_cast_1597_inst flow-through 
    process(type_cast_1597_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:type_cast_1597_inst:flowthrough inputs: " & " tmp1_1594 = "& Convert_SLV_To_Hex_String(tmp1_1594) & " outputs:" & " type_cast_1597_wire= "  & Convert_SLV_To_Hex_String(type_cast_1597_wire));
      --
    end process; 
    -- unary operator type_cast_1597_inst
    process(tmp1_1594) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp1_1594, tmp_var);
      type_cast_1597_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator ptr_deref_1539_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1539_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1539_load_0:started:   inputs: " & " ptr_deref_1539_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1539_word_address_0));
          --
        end if; 
        if ptr_deref_1539_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1539_load_0:finished:  outputs: " & " ptr_deref_1539_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1539_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_1469_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1469_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1469_load_0:started:   inputs: " & " ptr_deref_1469_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1469_word_address_0));
          --
        end if; 
        if ptr_deref_1469_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1469_load_0:finished:  outputs: " & " ptr_deref_1469_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1469_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : ptr_deref_1539_load_0 ptr_deref_1469_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1539_load_0_req_0,
        ptr_deref_1539_load_0_ack_0,
        ptr_deref_1539_load_0_req_1,
        ptr_deref_1539_load_0_ack_1,
        "ptr_deref_1539_load_0",
        "memory_space_3" ,
        ptr_deref_1539_data_0,
        ptr_deref_1539_word_address_0,
        "ptr_deref_1539_data_0",
        "ptr_deref_1539_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1469_load_0_req_0,
        ptr_deref_1469_load_0_ack_0,
        ptr_deref_1469_load_0_req_1,
        ptr_deref_1469_load_0_ack_1,
        "ptr_deref_1469_load_0",
        "memory_space_3" ,
        ptr_deref_1469_data_0,
        ptr_deref_1469_word_address_0,
        "ptr_deref_1469_data_0",
        "ptr_deref_1469_word_address_0" -- 
      );
      reqL_unguarded(1) <= ptr_deref_1539_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1469_load_0_req_0;
      ptr_deref_1539_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1469_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1539_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1469_load_0_req_1;
      ptr_deref_1539_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1469_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1539_word_address_0 & ptr_deref_1469_word_address_0;
      ptr_deref_1539_data_0 <= data_out(63 downto 32);
      ptr_deref_1469_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator ptr_deref_1638_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_1638_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1638_load_0:started:   inputs: " & " ptr_deref_1638_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_1638_word_address_0));
          --
        end if; 
        if ptr_deref_1638_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:ptr_deref_1638_load_0:finished:  outputs: " & " ptr_deref_1638_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_1638_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (1) : ptr_deref_1638_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1638_load_0_req_0,
        ptr_deref_1638_load_0_ack_0,
        ptr_deref_1638_load_0_req_1,
        ptr_deref_1638_load_0_ack_1,
        "ptr_deref_1638_load_0",
        "memory_space_0" ,
        ptr_deref_1638_data_0,
        ptr_deref_1638_word_address_0,
        "ptr_deref_1638_data_0",
        "ptr_deref_1638_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_1638_load_0_req_0;
      ptr_deref_1638_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1638_load_0_req_1;
      ptr_deref_1638_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1638_word_address_0;
      ptr_deref_1638_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- logger for split-operator WPIPE_maxpool_output_pipe_1677_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_maxpool_output_pipe_1677_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:WPIPE_maxpool_output_pipe_1677_inst:started:   PipeWrite to maxpool_output_pipe inputs: " & " conv35_1663 = "& Convert_SLV_To_Hex_String(conv35_1663));
          --
        end if; 
        if WPIPE_maxpool_output_pipe_1677_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:WPIPE_maxpool_output_pipe_1677_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator WPIPE_maxpool_output_pipe_1680_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_maxpool_output_pipe_1680_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:WPIPE_maxpool_output_pipe_1680_inst:started:   PipeWrite to maxpool_output_pipe inputs: " & " conv29_1653 = "& Convert_SLV_To_Hex_String(conv29_1653));
          --
        end if; 
        if WPIPE_maxpool_output_pipe_1680_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:WPIPE_maxpool_output_pipe_1680_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator WPIPE_maxpool_output_pipe_1683_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_maxpool_output_pipe_1683_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:WPIPE_maxpool_output_pipe_1683_inst:started:   PipeWrite to maxpool_output_pipe inputs: " & " conv23_1643 = "& Convert_SLV_To_Hex_String(conv23_1643));
          --
        end if; 
        if WPIPE_maxpool_output_pipe_1683_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:WPIPE_maxpool_output_pipe_1683_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator WPIPE_maxpool_output_pipe_1674_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_maxpool_output_pipe_1674_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:WPIPE_maxpool_output_pipe_1674_inst:started:   PipeWrite to maxpool_output_pipe inputs: " & " conv41_1673 = "& Convert_SLV_To_Hex_String(conv41_1673));
          --
        end if; 
        if WPIPE_maxpool_output_pipe_1674_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:sendB:DP:WPIPE_maxpool_output_pipe_1674_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1677_inst WPIPE_maxpool_output_pipe_1680_inst WPIPE_maxpool_output_pipe_1683_inst WPIPE_maxpool_output_pipe_1674_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1677_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1680_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1683_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1674_inst_req_0;
      WPIPE_maxpool_output_pipe_1677_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1680_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1683_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1674_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1677_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1680_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1683_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1674_inst_req_1;
      WPIPE_maxpool_output_pipe_1677_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1680_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1683_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1674_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      data_in <= conv35_1663 & conv29_1653 & conv23_1643 & conv41_1673;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(8 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(8 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    fill_T_call_reqs : out  std_logic_vector(0 downto 0);
    fill_T_call_acks : in   std_logic_vector(0 downto 0);
    fill_T_call_data : out  std_logic_vector(63 downto 0);
    fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
    fill_T_return_reqs : out  std_logic_vector(0 downto 0);
    fill_T_return_acks : in   std_logic_vector(0 downto 0);
    fill_T_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal testConfigure_CP_279_start: Boolean;
  signal testConfigure_CP_279_symbol: Boolean;
  -- volatile/operator module components. 
  component fill_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal if_stmt_299_branch_req_0 : boolean;
  signal call_stmt_373_call_req_1 : boolean;
  signal ptr_deref_281_load_2_ack_0 : boolean;
  signal ptr_deref_281_addr_1_req_1 : boolean;
  signal ptr_deref_212_addr_3_ack_1 : boolean;
  signal ptr_deref_281_load_2_req_0 : boolean;
  signal ptr_deref_212_addr_3_req_1 : boolean;
  signal if_stmt_219_branch_ack_0 : boolean;
  signal ptr_deref_281_addr_0_ack_0 : boolean;
  signal if_stmt_219_branch_ack_1 : boolean;
  signal ptr_deref_281_load_1_ack_0 : boolean;
  signal addr_of_277_final_reg_ack_1 : boolean;
  signal ptr_deref_281_load_1_req_0 : boolean;
  signal ptr_deref_281_load_0_ack_1 : boolean;
  signal array_obj_ref_276_index_offset_ack_1 : boolean;
  signal addr_of_277_final_reg_req_1 : boolean;
  signal array_obj_ref_276_index_offset_req_1 : boolean;
  signal ptr_deref_281_addr_1_ack_0 : boolean;
  signal ptr_deref_212_addr_3_ack_0 : boolean;
  signal ptr_deref_281_addr_1_req_0 : boolean;
  signal ptr_deref_281_load_0_ack_0 : boolean;
  signal ptr_deref_212_addr_3_req_0 : boolean;
  signal if_stmt_385_branch_ack_1 : boolean;
  signal if_stmt_385_branch_ack_0 : boolean;
  signal if_stmt_325_branch_ack_0 : boolean;
  signal ptr_deref_281_load_3_ack_1 : boolean;
  signal ptr_deref_281_addr_0_req_1 : boolean;
  signal ptr_deref_281_addr_0_req_0 : boolean;
  signal array_obj_ref_276_index_offset_ack_0 : boolean;
  signal array_obj_ref_276_index_offset_req_0 : boolean;
  signal ptr_deref_281_load_0_req_0 : boolean;
  signal if_stmt_219_branch_req_0 : boolean;
  signal ptr_deref_281_addr_0_ack_1 : boolean;
  signal ptr_deref_212_load_3_ack_0 : boolean;
  signal ptr_deref_212_load_3_req_0 : boolean;
  signal ptr_deref_281_load_3_ack_0 : boolean;
  signal ptr_deref_281_load_2_ack_1 : boolean;
  signal if_stmt_325_branch_ack_1 : boolean;
  signal ptr_deref_281_load_0_req_1 : boolean;
  signal if_stmt_299_branch_ack_1 : boolean;
  signal type_cast_341_inst_req_0 : boolean;
  signal type_cast_341_inst_ack_0 : boolean;
  signal if_stmt_325_branch_req_0 : boolean;
  signal type_cast_341_inst_req_1 : boolean;
  signal type_cast_341_inst_ack_1 : boolean;
  signal ptr_deref_281_load_1_ack_1 : boolean;
  signal if_stmt_385_branch_req_0 : boolean;
  signal ptr_deref_281_load_1_req_1 : boolean;
  signal array_obj_ref_276_index_1_scale_req_0 : boolean;
  signal if_stmt_137_branch_req_0 : boolean;
  signal if_stmt_137_branch_ack_1 : boolean;
  signal if_stmt_137_branch_ack_0 : boolean;
  signal call_stmt_373_call_req_0 : boolean;
  signal call_stmt_373_call_ack_0 : boolean;
  signal call_stmt_373_call_ack_1 : boolean;
  signal ptr_deref_212_load_2_ack_0 : boolean;
  signal ptr_deref_281_load_2_req_1 : boolean;
  signal if_stmt_299_branch_ack_0 : boolean;
  signal ptr_deref_212_addr_2_ack_1 : boolean;
  signal ptr_deref_281_load_3_req_1 : boolean;
  signal ptr_deref_212_load_2_req_0 : boolean;
  signal ptr_deref_212_load_1_ack_0 : boolean;
  signal addr_of_277_final_reg_ack_0 : boolean;
  signal ptr_deref_281_load_3_req_0 : boolean;
  signal ptr_deref_212_load_1_req_0 : boolean;
  signal ptr_deref_87_addr_0_req_0 : boolean;
  signal ptr_deref_87_addr_0_ack_0 : boolean;
  signal ptr_deref_212_addr_2_req_1 : boolean;
  signal ptr_deref_87_addr_0_req_1 : boolean;
  signal ptr_deref_87_addr_0_ack_1 : boolean;
  signal ptr_deref_87_addr_1_req_0 : boolean;
  signal ptr_deref_87_addr_1_ack_0 : boolean;
  signal ptr_deref_87_addr_1_req_1 : boolean;
  signal ptr_deref_87_addr_1_ack_1 : boolean;
  signal ptr_deref_87_addr_2_req_0 : boolean;
  signal ptr_deref_87_addr_2_ack_0 : boolean;
  signal ptr_deref_87_addr_2_req_1 : boolean;
  signal ptr_deref_87_addr_2_ack_1 : boolean;
  signal ptr_deref_87_addr_3_req_0 : boolean;
  signal ptr_deref_87_addr_3_ack_0 : boolean;
  signal ptr_deref_281_addr_3_ack_1 : boolean;
  signal ptr_deref_87_addr_3_req_1 : boolean;
  signal ptr_deref_87_addr_3_ack_1 : boolean;
  signal ptr_deref_281_addr_3_req_1 : boolean;
  signal ptr_deref_87_store_0_req_0 : boolean;
  signal ptr_deref_87_store_0_ack_0 : boolean;
  signal ptr_deref_87_store_1_req_0 : boolean;
  signal ptr_deref_87_store_1_ack_0 : boolean;
  signal ptr_deref_212_addr_2_ack_0 : boolean;
  signal ptr_deref_87_store_2_req_0 : boolean;
  signal ptr_deref_87_store_2_ack_0 : boolean;
  signal ptr_deref_87_store_3_req_0 : boolean;
  signal ptr_deref_87_store_3_ack_0 : boolean;
  signal ptr_deref_281_addr_3_ack_0 : boolean;
  signal ptr_deref_87_store_0_req_1 : boolean;
  signal ptr_deref_87_store_0_ack_1 : boolean;
  signal ptr_deref_281_addr_3_req_0 : boolean;
  signal ptr_deref_87_store_1_req_1 : boolean;
  signal ptr_deref_87_store_1_ack_1 : boolean;
  signal ptr_deref_212_addr_2_req_0 : boolean;
  signal ptr_deref_87_store_2_req_1 : boolean;
  signal ptr_deref_87_store_2_ack_1 : boolean;
  signal ptr_deref_87_store_3_req_1 : boolean;
  signal ptr_deref_87_store_3_ack_1 : boolean;
  signal addr_of_277_final_reg_req_0 : boolean;
  signal ptr_deref_212_load_0_ack_0 : boolean;
  signal ptr_deref_212_load_0_req_0 : boolean;
  signal ptr_deref_98_store_0_req_0 : boolean;
  signal ptr_deref_98_store_0_ack_0 : boolean;
  signal ptr_deref_98_store_0_req_1 : boolean;
  signal ptr_deref_98_store_0_ack_1 : boolean;
  signal array_obj_ref_276_index_1_scale_ack_1 : boolean;
  signal array_obj_ref_276_index_1_scale_req_1 : boolean;
  signal ptr_deref_109_addr_0_req_0 : boolean;
  signal ptr_deref_109_addr_0_ack_0 : boolean;
  signal ptr_deref_281_addr_2_ack_1 : boolean;
  signal ptr_deref_109_addr_0_req_1 : boolean;
  signal ptr_deref_109_addr_0_ack_1 : boolean;
  signal ptr_deref_212_addr_1_ack_1 : boolean;
  signal ptr_deref_281_addr_2_req_1 : boolean;
  signal ptr_deref_109_addr_1_req_0 : boolean;
  signal ptr_deref_109_addr_1_ack_0 : boolean;
  signal ptr_deref_212_addr_1_req_1 : boolean;
  signal ptr_deref_109_addr_1_req_1 : boolean;
  signal ptr_deref_109_addr_1_ack_1 : boolean;
  signal ptr_deref_109_addr_2_req_0 : boolean;
  signal ptr_deref_109_addr_2_ack_0 : boolean;
  signal ptr_deref_109_addr_2_req_1 : boolean;
  signal ptr_deref_109_addr_2_ack_1 : boolean;
  signal ptr_deref_212_addr_1_ack_0 : boolean;
  signal ptr_deref_109_addr_3_req_0 : boolean;
  signal ptr_deref_109_addr_3_ack_0 : boolean;
  signal ptr_deref_212_addr_1_req_0 : boolean;
  signal ptr_deref_281_addr_2_ack_0 : boolean;
  signal ptr_deref_109_addr_3_req_1 : boolean;
  signal type_cast_240_inst_ack_1 : boolean;
  signal ptr_deref_109_addr_3_ack_1 : boolean;
  signal type_cast_240_inst_req_1 : boolean;
  signal ptr_deref_281_addr_2_req_0 : boolean;
  signal ptr_deref_109_store_0_req_0 : boolean;
  signal ptr_deref_109_store_0_ack_0 : boolean;
  signal ptr_deref_109_store_1_req_0 : boolean;
  signal ptr_deref_109_store_1_ack_0 : boolean;
  signal ptr_deref_109_store_2_req_0 : boolean;
  signal ptr_deref_109_store_2_ack_0 : boolean;
  signal ptr_deref_195_store_0_ack_1 : boolean;
  signal ptr_deref_109_store_3_req_0 : boolean;
  signal ptr_deref_109_store_3_ack_0 : boolean;
  signal ptr_deref_195_store_0_req_1 : boolean;
  signal ptr_deref_109_store_0_req_1 : boolean;
  signal type_cast_240_inst_ack_0 : boolean;
  signal ptr_deref_109_store_0_ack_1 : boolean;
  signal ptr_deref_109_store_1_req_1 : boolean;
  signal ptr_deref_109_store_1_ack_1 : boolean;
  signal ptr_deref_212_addr_0_ack_1 : boolean;
  signal ptr_deref_109_store_2_req_1 : boolean;
  signal type_cast_240_inst_req_0 : boolean;
  signal ptr_deref_109_store_2_ack_1 : boolean;
  signal ptr_deref_109_store_3_req_1 : boolean;
  signal ptr_deref_212_addr_0_req_1 : boolean;
  signal ptr_deref_109_store_3_ack_1 : boolean;
  signal array_obj_ref_276_index_1_scale_ack_0 : boolean;
  signal ptr_deref_212_addr_0_ack_0 : boolean;
  signal ptr_deref_212_load_3_ack_1 : boolean;
  signal ptr_deref_212_load_3_req_1 : boolean;
  signal ptr_deref_212_addr_0_req_0 : boolean;
  signal ptr_deref_212_load_2_ack_1 : boolean;
  signal ptr_deref_212_load_2_req_1 : boolean;
  signal ptr_deref_120_store_0_req_0 : boolean;
  signal ptr_deref_120_store_0_ack_0 : boolean;
  signal ptr_deref_281_addr_1_ack_1 : boolean;
  signal ptr_deref_120_store_0_req_1 : boolean;
  signal ptr_deref_212_load_1_ack_1 : boolean;
  signal ptr_deref_120_store_0_ack_1 : boolean;
  signal ptr_deref_212_load_1_req_1 : boolean;
  signal ptr_deref_212_load_0_ack_1 : boolean;
  signal ptr_deref_212_load_0_req_1 : boolean;
  signal type_cast_160_inst_req_0 : boolean;
  signal type_cast_160_inst_ack_0 : boolean;
  signal type_cast_160_inst_req_1 : boolean;
  signal type_cast_160_inst_ack_1 : boolean;
  signal array_obj_ref_166_index_offset_req_0 : boolean;
  signal array_obj_ref_166_index_offset_ack_0 : boolean;
  signal array_obj_ref_166_index_offset_req_1 : boolean;
  signal array_obj_ref_166_index_offset_ack_1 : boolean;
  signal addr_of_167_final_reg_req_0 : boolean;
  signal addr_of_167_final_reg_ack_0 : boolean;
  signal addr_of_167_final_reg_req_1 : boolean;
  signal addr_of_167_final_reg_ack_1 : boolean;
  signal array_obj_ref_173_index_1_scale_req_0 : boolean;
  signal array_obj_ref_173_index_1_scale_ack_0 : boolean;
  signal array_obj_ref_173_index_1_scale_req_1 : boolean;
  signal array_obj_ref_173_index_1_scale_ack_1 : boolean;
  signal array_obj_ref_173_index_offset_req_0 : boolean;
  signal array_obj_ref_173_index_offset_ack_0 : boolean;
  signal array_obj_ref_173_index_offset_req_1 : boolean;
  signal array_obj_ref_173_index_offset_ack_1 : boolean;
  signal addr_of_174_final_reg_req_0 : boolean;
  signal addr_of_174_final_reg_ack_0 : boolean;
  signal addr_of_174_final_reg_req_1 : boolean;
  signal addr_of_174_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_177_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_177_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_177_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_177_inst_ack_1 : boolean;
  signal type_cast_181_inst_req_0 : boolean;
  signal type_cast_181_inst_ack_0 : boolean;
  signal type_cast_181_inst_req_1 : boolean;
  signal type_cast_181_inst_ack_1 : boolean;
  signal ptr_deref_184_addr_0_req_0 : boolean;
  signal ptr_deref_184_addr_0_ack_0 : boolean;
  signal ptr_deref_184_addr_0_req_1 : boolean;
  signal ptr_deref_184_addr_0_ack_1 : boolean;
  signal ptr_deref_184_addr_1_req_0 : boolean;
  signal ptr_deref_184_addr_1_ack_0 : boolean;
  signal ptr_deref_184_addr_1_req_1 : boolean;
  signal ptr_deref_184_addr_1_ack_1 : boolean;
  signal ptr_deref_184_addr_2_req_0 : boolean;
  signal ptr_deref_184_addr_2_ack_0 : boolean;
  signal ptr_deref_184_addr_2_req_1 : boolean;
  signal ptr_deref_184_addr_2_ack_1 : boolean;
  signal ptr_deref_184_addr_3_req_0 : boolean;
  signal ptr_deref_184_addr_3_ack_0 : boolean;
  signal ptr_deref_184_addr_3_req_1 : boolean;
  signal ptr_deref_184_addr_3_ack_1 : boolean;
  signal ptr_deref_184_store_0_req_0 : boolean;
  signal ptr_deref_184_store_0_ack_0 : boolean;
  signal ptr_deref_184_store_1_req_0 : boolean;
  signal ptr_deref_184_store_1_ack_0 : boolean;
  signal ptr_deref_184_store_2_req_0 : boolean;
  signal ptr_deref_184_store_2_ack_0 : boolean;
  signal ptr_deref_184_store_3_req_0 : boolean;
  signal ptr_deref_184_store_3_ack_0 : boolean;
  signal ptr_deref_184_store_0_req_1 : boolean;
  signal ptr_deref_184_store_0_ack_1 : boolean;
  signal ptr_deref_184_store_1_req_1 : boolean;
  signal ptr_deref_184_store_1_ack_1 : boolean;
  signal ptr_deref_184_store_2_req_1 : boolean;
  signal ptr_deref_184_store_2_ack_1 : boolean;
  signal ptr_deref_184_store_3_req_1 : boolean;
  signal ptr_deref_184_store_3_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_188_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_188_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_188_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_188_inst_ack_1 : boolean;
  signal type_cast_192_inst_req_0 : boolean;
  signal type_cast_192_inst_ack_0 : boolean;
  signal type_cast_192_inst_req_1 : boolean;
  signal type_cast_192_inst_ack_1 : boolean;
  signal ptr_deref_195_store_0_req_0 : boolean;
  signal ptr_deref_195_store_0_ack_0 : boolean;
  signal type_cast_129_inst_req_0 : boolean;
  signal type_cast_129_inst_ack_0 : boolean;
  signal type_cast_129_inst_req_1 : boolean;
  signal type_cast_129_inst_ack_1 : boolean;
  signal phi_stmt_126_req_0 : boolean;
  signal phi_stmt_126_ack_0 : boolean;
  signal phi_stmt_144_req_0 : boolean;
  signal type_cast_150_inst_req_0 : boolean;
  signal type_cast_150_inst_ack_0 : boolean;
  signal type_cast_150_inst_req_1 : boolean;
  signal type_cast_150_inst_ack_1 : boolean;
  signal phi_stmt_144_req_1 : boolean;
  signal phi_stmt_144_ack_0 : boolean;
  signal phi_stmt_257_req_0 : boolean;
  signal phi_stmt_264_req_0 : boolean;
  signal type_cast_263_inst_req_0 : boolean;
  signal type_cast_263_inst_ack_0 : boolean;
  signal type_cast_263_inst_req_1 : boolean;
  signal type_cast_263_inst_ack_1 : boolean;
  signal phi_stmt_257_req_1 : boolean;
  signal type_cast_270_inst_req_0 : boolean;
  signal type_cast_270_inst_ack_0 : boolean;
  signal type_cast_270_inst_req_1 : boolean;
  signal type_cast_270_inst_ack_1 : boolean;
  signal phi_stmt_264_req_1 : boolean;
  signal phi_stmt_257_ack_0 : boolean;
  signal phi_stmt_264_ack_0 : boolean;
  signal type_cast_313_inst_req_0 : boolean;
  signal type_cast_313_inst_ack_0 : boolean;
  signal type_cast_313_inst_req_1 : boolean;
  signal type_cast_313_inst_ack_1 : boolean;
  signal phi_stmt_310_req_0 : boolean;
  signal type_cast_309_inst_req_0 : boolean;
  signal type_cast_309_inst_ack_0 : boolean;
  signal type_cast_309_inst_req_1 : boolean;
  signal type_cast_309_inst_ack_1 : boolean;
  signal phi_stmt_306_req_0 : boolean;
  signal type_cast_317_inst_req_0 : boolean;
  signal type_cast_317_inst_ack_0 : boolean;
  signal type_cast_317_inst_req_1 : boolean;
  signal type_cast_317_inst_ack_1 : boolean;
  signal phi_stmt_314_req_0 : boolean;
  signal phi_stmt_306_ack_0 : boolean;
  signal phi_stmt_310_ack_0 : boolean;
  signal phi_stmt_314_ack_0 : boolean;
  signal phi_stmt_364_req_0 : boolean;
  signal type_cast_370_inst_req_0 : boolean;
  signal type_cast_370_inst_ack_0 : boolean;
  signal type_cast_370_inst_req_1 : boolean;
  signal type_cast_370_inst_ack_1 : boolean;
  signal phi_stmt_364_req_1 : boolean;
  signal phi_stmt_364_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_279_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_279_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_279_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_279_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,testConfigure_CP_279_start,"testConfigure cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,testConfigure_CP_279_symbol, "testConfigure cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_279: Block -- control-path 
    signal testConfigure_CP_279_elements: BooleanArray(207 downto 0);
    -- 
  begin -- 
    testConfigure_CP_279_elements(0) <= testConfigure_CP_279_start;
    testConfigure_CP_279_symbol <= testConfigure_CP_279_elements(207);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	26 
    -- CP-element group 0: 	47 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	30 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	35 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	42 
    -- CP-element group 0: 	43 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	18 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	23 
    -- CP-element group 0:  members (136) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_79/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/branch_block_stmt_79__entry__
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123__entry__
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_update_start_
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_sample_start
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_update_start
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_0_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_0_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_0_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_0_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_1_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_1_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_1_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_1_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_2_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_2_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_2_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_2_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_3_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_3_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_3_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_3_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_1/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_2/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_2/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_3/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_3/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_update_start_
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_update_start_
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_sample_start
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_update_start
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_0_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_0_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_0_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_0_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_1_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_1_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_1_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_1_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_2_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_2_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_2_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_2_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_3_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_3_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_3_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_3_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_1/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_2/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_2/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_3/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_3/cr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_update_start_
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/ptr_deref_120_Split/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/ptr_deref_120_Split/$exit
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/ptr_deref_120_Split/split_req
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/ptr_deref_120_Split/split_ack
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_3_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_98_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_3_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_120_store_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_120_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_addr_0_req_0); -- 
    cr_366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_addr_0_req_1); -- 
    rr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_addr_1_req_0); -- 
    cr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_addr_1_req_1); -- 
    rr_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_addr_2_req_0); -- 
    cr_386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_addr_2_req_1); -- 
    rr_391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_addr_3_req_0); -- 
    cr_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_addr_3_req_1); -- 
    cr_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_store_0_req_1); -- 
    cr_443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_store_1_req_1); -- 
    cr_448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_store_2_req_1); -- 
    cr_453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_87_store_3_req_1); -- 
    cr_503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_98_store_0_req_1); -- 
    rr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_addr_0_req_0); -- 
    cr_535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_addr_0_req_1); -- 
    rr_540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_addr_1_req_0); -- 
    cr_545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_addr_1_req_1); -- 
    rr_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_addr_2_req_0); -- 
    cr_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_addr_2_req_1); -- 
    rr_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_addr_3_req_0); -- 
    cr_565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_addr_3_req_1); -- 
    cr_607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_store_0_req_1); -- 
    cr_612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_store_1_req_1); -- 
    cr_617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_store_2_req_1); -- 
    cr_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_109_store_3_req_1); -- 
    rr_661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_120_store_0_req_0); -- 
    cr_672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(0), ack => ptr_deref_120_store_0_req_1); -- 
    -- CP-element group 1:  merge  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	200 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	155 
    -- CP-element group 1: 	156 
    -- CP-element group 1:  members (13) 
      -- CP-element group 1: 	 branch_block_stmt_79/if_stmt_325_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_79/if_stmt_325_else_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_79/R_cmp3445_326_place
      -- CP-element group 1: 	 branch_block_stmt_79/assign_stmt_324/$entry
      -- CP-element group 1: 	 branch_block_stmt_79/assign_stmt_324/$exit
      -- CP-element group 1: 	 branch_block_stmt_79/if_stmt_325_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_79/if_stmt_325_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_79/if_stmt_325_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_79/if_stmt_325_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_79/merge_stmt_305__exit__
      -- CP-element group 1: 	 branch_block_stmt_79/assign_stmt_324__entry__
      -- CP-element group 1: 	 branch_block_stmt_79/assign_stmt_324__exit__
      -- CP-element group 1: 	 branch_block_stmt_79/if_stmt_325__entry__
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_325_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_1403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(1), ack => if_stmt_325_branch_req_0); -- 
    testConfigure_CP_279_elements(1) <= testConfigure_CP_279_elements(200);
    -- CP-element group 2:  join  fork  transition  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: 	4 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2:  members (15) 
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/ptr_deref_87_Split/$entry
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/ptr_deref_87_Split/$exit
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/ptr_deref_87_Split/split_req
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/ptr_deref_87_Split/split_ack
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_1/$entry
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_1/rr
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_2/$entry
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_2/rr
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_3/$entry
      -- CP-element group 2: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_3/rr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_3_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(2), ack => ptr_deref_87_store_0_req_0); -- 
    rr_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(2), ack => ptr_deref_87_store_1_req_0); -- 
    rr_422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(2), ack => ptr_deref_87_store_2_req_0); -- 
    rr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(2), ack => ptr_deref_87_store_3_req_0); -- 
    testConfigure_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(0) & testConfigure_CP_279_elements(4);
      gj_testConfigure_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	5 
    -- CP-element group 3: 	7 
    -- CP-element group 3: 	9 
    -- CP-element group 3: 	11 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	51 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_sample_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(5) & testConfigure_CP_279_elements(7) & testConfigure_CP_279_elements(9) & testConfigure_CP_279_elements(11);
      gj_testConfigure_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	8 
    -- CP-element group 4: 	10 
    -- CP-element group 4: 	12 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	2 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_address_calculated
      -- CP-element group 4: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_update_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(6) & testConfigure_CP_279_elements(8) & testConfigure_CP_279_elements(10) & testConfigure_CP_279_elements(12);
      gj_testConfigure_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	3 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_0_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_0_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_addr_0_ack_0, ack => testConfigure_CP_279_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	4 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_0_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_0_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_addr_0_ack_1, ack => testConfigure_CP_279_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	3 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_1_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_1_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_addr_1_ack_0, ack => testConfigure_CP_279_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	4 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_1_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_1_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_addr_1_ack_1, ack => testConfigure_CP_279_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	3 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_2_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_2_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_addr_2_ack_0, ack => testConfigure_CP_279_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	4 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_2_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_2_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_addr_2_ack_1, ack => testConfigure_CP_279_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	3 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_3_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_3_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_addr_3_ack_0, ack => testConfigure_CP_279_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	4 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_3_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_word_addrgen_3_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_addr_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_addr_3_ack_1, ack => testConfigure_CP_279_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	17 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_store_0_ack_0, ack => testConfigure_CP_279_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_1/$exit
      -- CP-element group 14: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_1/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_store_1_ack_0, ack => testConfigure_CP_279_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_2/$exit
      -- CP-element group 15: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_2/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_store_2_ack_0, ack => testConfigure_CP_279_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_3/$exit
      -- CP-element group 16: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/word_3/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_store_3_ack_0, ack => testConfigure_CP_279_elements(16)); -- 
    -- CP-element group 17:  join  transition  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	13 
    -- CP-element group 17: 	14 
    -- CP-element group 17: 	15 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	49 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(13) & testConfigure_CP_279_elements(14) & testConfigure_CP_279_elements(15) & testConfigure_CP_279_elements(16);
      gj_testConfigure_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	0 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_store_0_ack_1, ack => testConfigure_CP_279_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_1/$exit
      -- CP-element group 19: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_1/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_store_1_ack_1, ack => testConfigure_CP_279_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_2/$exit
      -- CP-element group 20: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_2/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_store_2_ack_1, ack => testConfigure_CP_279_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_3/$exit
      -- CP-element group 21: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/word_3/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_87_store_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_87_store_3_ack_1, ack => testConfigure_CP_279_elements(21)); -- 
    -- CP-element group 22:  join  transition  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: 	19 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	51 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_Update/word_access_complete/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(18) & testConfigure_CP_279_elements(19) & testConfigure_CP_279_elements(20) & testConfigure_CP_279_elements(21);
      gj_testConfigure_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: 	49 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/ptr_deref_98_Split/$entry
      -- CP-element group 23: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/ptr_deref_98_Split/$exit
      -- CP-element group 23: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/ptr_deref_98_Split/split_req
      -- CP-element group 23: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/ptr_deref_98_Split/split_ack
      -- CP-element group 23: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/word_access_start/$entry
      -- CP-element group 23: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_98_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(23), ack => ptr_deref_98_store_0_req_0); -- 
    testConfigure_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(0) & testConfigure_CP_279_elements(49);
      gj_testConfigure_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	50 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/word_access_start/$exit
      -- CP-element group 24: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_98_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_98_store_0_ack_0, ack => testConfigure_CP_279_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	51 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Update/word_access_complete/$exit
      -- CP-element group 25: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_98_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_98_store_0_ack_1, ack => testConfigure_CP_279_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: 	28 
    -- CP-element group 26: 	50 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	37 
    -- CP-element group 26: 	38 
    -- CP-element group 26: 	39 
    -- CP-element group 26: 	40 
    -- CP-element group 26:  members (15) 
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/ptr_deref_109_Split/$entry
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/ptr_deref_109_Split/$exit
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/ptr_deref_109_Split/split_req
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/ptr_deref_109_Split/split_ack
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/$entry
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_0/$entry
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_0/rr
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_1/$entry
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_1/rr
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_2/$entry
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_2/rr
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_3/$entry
      -- CP-element group 26: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_3/rr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_3_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(26), ack => ptr_deref_109_store_0_req_0); -- 
    rr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(26), ack => ptr_deref_109_store_1_req_0); -- 
    rr_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(26), ack => ptr_deref_109_store_2_req_0); -- 
    rr_596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(26), ack => ptr_deref_109_store_3_req_0); -- 
    testConfigure_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(0) & testConfigure_CP_279_elements(28) & testConfigure_CP_279_elements(50);
      gj_testConfigure_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: 	31 
    -- CP-element group 27: 	33 
    -- CP-element group 27: 	35 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	51 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_sample_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(27) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(29) & testConfigure_CP_279_elements(31) & testConfigure_CP_279_elements(33) & testConfigure_CP_279_elements(35);
      gj_testConfigure_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: 	32 
    -- CP-element group 28: 	34 
    -- CP-element group 28: 	36 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_address_calculated
      -- CP-element group 28: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_update_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(30) & testConfigure_CP_279_elements(32) & testConfigure_CP_279_elements(34) & testConfigure_CP_279_elements(36);
      gj_testConfigure_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_0_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_0_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_addr_0_ack_0, ack => testConfigure_CP_279_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	0 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_0_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_0_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_addr_0_ack_1, ack => testConfigure_CP_279_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	27 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_1_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_1_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_addr_1_ack_0, ack => testConfigure_CP_279_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	28 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_1_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_1_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_addr_1_ack_1, ack => testConfigure_CP_279_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	27 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_2_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_2_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_addr_2_ack_0, ack => testConfigure_CP_279_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	0 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	28 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_2_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_2_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_addr_2_ack_1, ack => testConfigure_CP_279_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	0 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	27 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_3_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_3_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_addr_3_ack_0, ack => testConfigure_CP_279_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	28 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_3_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_word_addrgen_3_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_addr_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_addr_3_ack_1, ack => testConfigure_CP_279_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	26 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	41 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_store_0_ack_0, ack => testConfigure_CP_279_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	26 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_1/$exit
      -- CP-element group 38: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_1/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_store_1_ack_0, ack => testConfigure_CP_279_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	26 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_2/$exit
      -- CP-element group 39: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_2/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_store_2_ack_0, ack => testConfigure_CP_279_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	26 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_3/$exit
      -- CP-element group 40: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/word_3/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_store_3_ack_0, ack => testConfigure_CP_279_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	37 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(41) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(37) & testConfigure_CP_279_elements(38) & testConfigure_CP_279_elements(39) & testConfigure_CP_279_elements(40);
      gj_testConfigure_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	0 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	46 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_store_0_ack_1, ack => testConfigure_CP_279_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	0 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_1/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_store_1_ack_1, ack => testConfigure_CP_279_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_2/$exit
      -- CP-element group 44: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_2/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_store_2_ack_1, ack => testConfigure_CP_279_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_3/$exit
      -- CP-element group 45: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/word_3/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_109_store_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_109_store_3_ack_1, ack => testConfigure_CP_279_elements(45)); -- 
    -- CP-element group 46:  join  transition  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	42 
    -- CP-element group 46: 	43 
    -- CP-element group 46: 	44 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	51 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_109_Update/word_access_complete/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(42) & testConfigure_CP_279_elements(43) & testConfigure_CP_279_elements(44) & testConfigure_CP_279_elements(45);
      gj_testConfigure_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	0 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/word_access_start/$exit
      -- CP-element group 47: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/word_access_start/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_120_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_120_store_0_ack_0, ack => testConfigure_CP_279_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	51 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Update/word_access_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Update/word_access_complete/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_120_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_120_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_120_store_0_ack_1, ack => testConfigure_CP_279_elements(48)); -- 
    -- CP-element group 49:  transition  delay-element  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	23 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_87_ptr_deref_98_delay
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(49) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group testConfigure_CP_279_elements(49) is a control-delay.
    cp_element_49_delay: control_delay_element  generic map(name => " 49_delay", delay_value => 1)  port map(req => testConfigure_CP_279_elements(17), ack => testConfigure_CP_279_elements(49), clk => clk, reset =>reset);
    -- CP-element group 50:  transition  delay-element  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	24 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	26 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/ptr_deref_98_ptr_deref_109_delay
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(50) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group testConfigure_CP_279_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => testConfigure_CP_279_elements(24), ack => testConfigure_CP_279_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  transition  place  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	46 
    -- CP-element group 51: 	25 
    -- CP-element group 51: 	27 
    -- CP-element group 51: 	48 
    -- CP-element group 51: 	3 
    -- CP-element group 51: 	22 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	167 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123__exit__
      -- CP-element group 51: 	 branch_block_stmt_79/bbx_xnph55_forx_xbody
      -- CP-element group 51: 	 branch_block_stmt_79/assign_stmt_85_to_assign_stmt_123/$exit
      -- CP-element group 51: 	 branch_block_stmt_79/bbx_xnph55_forx_xbody_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_79/bbx_xnph55_forx_xbody_PhiReq/phi_stmt_144/$entry
      -- CP-element group 51: 	 branch_block_stmt_79/bbx_xnph55_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(46) & testConfigure_CP_279_elements(25) & testConfigure_CP_279_elements(27) & testConfigure_CP_279_elements(48) & testConfigure_CP_279_elements(3) & testConfigure_CP_279_elements(22);
      gj_testConfigure_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  place  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	166 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	207 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_79/if_stmt_137_if_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_79/if_stmt_137_if_link/if_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_79/forx_xcond13x_xpreheader_forx_xend42
      -- CP-element group 52: 	 branch_block_stmt_79/forx_xcond13x_xpreheader_forx_xend42_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_79/forx_xcond13x_xpreheader_forx_xend42_PhiReq/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_137_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_137_branch_ack_1, ack => testConfigure_CP_279_elements(52)); -- 
    -- CP-element group 53:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	166 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	123 
    -- CP-element group 53: 	124 
    -- CP-element group 53:  members (18) 
      -- CP-element group 53: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/$entry
      -- CP-element group 53: 	 branch_block_stmt_79/if_stmt_137_else_link/$exit
      -- CP-element group 53: 	 branch_block_stmt_79/if_stmt_137_else_link/else_choice_transition
      -- CP-element group 53: 	 branch_block_stmt_79/forx_xcond13x_xpreheader_bbx_xnph51
      -- CP-element group 53: 	 branch_block_stmt_79/merge_stmt_225__exit__
      -- CP-element group 53: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254__entry__
      -- CP-element group 53: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_Update/cr
      -- CP-element group 53: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_update_start_
      -- CP-element group 53: 	 branch_block_stmt_79/forx_xcond13x_xpreheader_bbx_xnph51_PhiReq/$entry
      -- CP-element group 53: 	 branch_block_stmt_79/forx_xcond13x_xpreheader_bbx_xnph51_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_79/merge_stmt_225_PhiReqMerge
      -- CP-element group 53: 	 branch_block_stmt_79/merge_stmt_225_PhiAck/$entry
      -- CP-element group 53: 	 branch_block_stmt_79/merge_stmt_225_PhiAck/$exit
      -- CP-element group 53: 	 branch_block_stmt_79/merge_stmt_225_PhiAck/dummy
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_137_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_240_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_240_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_137_branch_ack_0, ack => testConfigure_CP_279_elements(53)); -- 
    cr_1195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(53), ack => type_cast_240_inst_req_1); -- 
    rr_1190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(53), ack => type_cast_240_inst_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	172 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_160_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_160_inst_ack_0, ack => testConfigure_CP_279_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	172 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	120 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_160_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_160_inst_ack_1, ack => testConfigure_CP_279_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	172 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	120 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_final_index_sum_regn_sample_complete
      -- CP-element group 56: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_final_index_sum_regn_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_166_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_166_index_offset_ack_0, ack => testConfigure_CP_279_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	172 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (11) 
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_root_address_calculated
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_offset_calculated
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_final_index_sum_regn_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_final_index_sum_regn_Update/ack
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_base_plus_offset/$entry
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_base_plus_offset/$exit
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_base_plus_offset/sum_rename_req
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_base_plus_offset/sum_rename_ack
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_request/$entry
      -- CP-element group 57: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_request/req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_166_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_167_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_166_index_offset_ack_1, ack => testConfigure_CP_279_elements(57)); -- 
    req_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(57), ack => addr_of_167_final_reg_req_0); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_request/$exit
      -- CP-element group 58: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_request/ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_167_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_167_final_reg_ack_0, ack => testConfigure_CP_279_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	172 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	95 
    -- CP-element group 59:  members (19) 
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_complete/$exit
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_complete/ack
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_base_address_calculated
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_word_address_calculated
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_root_address_calculated
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_base_address_resized
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_base_addr_resize/$entry
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_base_addr_resize/$exit
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_base_addr_resize/base_resize_req
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_base_addr_resize/base_resize_ack
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_base_plus_offset/$entry
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_base_plus_offset/$exit
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_base_plus_offset/sum_rename_req
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_base_plus_offset/sum_rename_ack
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_word_addrgen/$entry
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_word_addrgen/$exit
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_word_addrgen/root_register_req
      -- CP-element group 59: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_167_final_reg_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_167_final_reg_ack_1, ack => testConfigure_CP_279_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	172 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	120 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_sample_complete
      -- CP-element group 60: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_173_index_1_scale_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_173_index_1_scale_ack_0, ack => testConfigure_CP_279_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	172 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scaled_1
      -- CP-element group 61: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_update_complete
      -- CP-element group 61: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_final_index_sum_regn_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_final_index_sum_regn_Sample/req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_173_index_1_scale_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_173_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_173_index_1_scale_ack_1, ack => testConfigure_CP_279_elements(61)); -- 
    req_794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(61), ack => array_obj_ref_173_index_offset_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	120 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_final_index_sum_regn_sample_complete
      -- CP-element group 62: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_final_index_sum_regn_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_173_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_173_index_offset_ack_0, ack => testConfigure_CP_279_elements(62)); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	172 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (11) 
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_root_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_offset_calculated
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_final_index_sum_regn_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_final_index_sum_regn_Update/ack
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_base_plus_offset/$entry
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_base_plus_offset/$exit
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_base_plus_offset/sum_rename_req
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_base_plus_offset/sum_rename_ack
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_request/$entry
      -- CP-element group 63: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_request/req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_173_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_174_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_173_index_offset_ack_1, ack => testConfigure_CP_279_elements(63)); -- 
    req_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(63), ack => addr_of_174_final_reg_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_request/$exit
      -- CP-element group 64: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_request/ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_174_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_174_final_reg_ack_0, ack => testConfigure_CP_279_elements(64)); -- 
    -- CP-element group 65:  fork  transition  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	172 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	70 
    -- CP-element group 65: 	73 
    -- CP-element group 65: 	75 
    -- CP-element group 65: 	77 
    -- CP-element group 65: 	79 
    -- CP-element group 65:  members (23) 
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_complete/ack
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_base_address_calculated
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_root_address_calculated
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_base_address_resized
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_base_addr_resize/$entry
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_base_addr_resize/$exit
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_base_addr_resize/base_resize_req
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_base_addr_resize/base_resize_ack
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_base_plus_offset/$entry
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_base_plus_offset/$exit
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_base_plus_offset/sum_rename_req
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_base_plus_offset/sum_rename_ack
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_sample_start
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_0_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_0_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_1_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_1_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_2_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_2_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_3_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_3_Sample/rr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_174_final_reg_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_3_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_174_final_reg_ack_1, ack => testConfigure_CP_279_elements(65)); -- 
    rr_869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(65), ack => ptr_deref_184_addr_0_req_0); -- 
    rr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(65), ack => ptr_deref_184_addr_1_req_0); -- 
    rr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(65), ack => ptr_deref_184_addr_2_req_0); -- 
    rr_899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(65), ack => ptr_deref_184_addr_3_req_0); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	172 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_update_start_
      -- CP-element group 66: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_Update/cr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:RPIPE_maxpool_input_pipe_177_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:RPIPE_maxpool_input_pipe_177_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_177_inst_ack_0, ack => testConfigure_CP_279_elements(66)); -- 
    cr_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(66), ack => RPIPE_maxpool_input_pipe_177_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	91 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_Sample/rr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:RPIPE_maxpool_input_pipe_177_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_181_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:RPIPE_maxpool_input_pipe_188_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_177_inst_ack_1, ack => testConfigure_CP_279_elements(67)); -- 
    rr_837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(67), ack => type_cast_181_inst_req_0); -- 
    rr_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(67), ack => RPIPE_maxpool_input_pipe_188_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_181_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_181_inst_ack_0, ack => testConfigure_CP_279_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	172 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_181_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_181_inst_ack_1, ack => testConfigure_CP_279_elements(69)); -- 
    -- CP-element group 70:  join  fork  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	65 
    -- CP-element group 70: 	69 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	81 
    -- CP-element group 70: 	82 
    -- CP-element group 70: 	83 
    -- CP-element group 70: 	84 
    -- CP-element group 70:  members (15) 
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/ptr_deref_184_Split/$entry
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/ptr_deref_184_Split/$exit
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/ptr_deref_184_Split/split_req
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/ptr_deref_184_Split/split_ack
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/$entry
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_0/$entry
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_0/rr
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_1/$entry
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_1/rr
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_2/$entry
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_2/rr
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_3/$entry
      -- CP-element group 70: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_3/rr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_3_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(70), ack => ptr_deref_184_store_0_req_0); -- 
    rr_925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(70), ack => ptr_deref_184_store_1_req_0); -- 
    rr_930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(70), ack => ptr_deref_184_store_2_req_0); -- 
    rr_935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(70), ack => ptr_deref_184_store_3_req_0); -- 
    testConfigure_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(65) & testConfigure_CP_279_elements(69) & testConfigure_CP_279_elements(72);
      gj_testConfigure_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	75 
    -- CP-element group 71: 	77 
    -- CP-element group 71: 	79 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	120 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_sample_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(71) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(73) & testConfigure_CP_279_elements(75) & testConfigure_CP_279_elements(77) & testConfigure_CP_279_elements(79);
      gj_testConfigure_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  join  transition  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: 	76 
    -- CP-element group 72: 	78 
    -- CP-element group 72: 	80 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_update_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(72) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(74) & testConfigure_CP_279_elements(76) & testConfigure_CP_279_elements(78) & testConfigure_CP_279_elements(80);
      gj_testConfigure_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	65 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_0_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_0_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_addr_0_ack_0, ack => testConfigure_CP_279_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	172 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	72 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_0_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_0_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_addr_0_ack_1, ack => testConfigure_CP_279_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	65 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	71 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_1_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_1_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_addr_1_ack_0, ack => testConfigure_CP_279_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	172 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	72 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_1_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_1_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_addr_1_ack_1, ack => testConfigure_CP_279_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	65 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	71 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_2_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_2_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_addr_2_ack_0, ack => testConfigure_CP_279_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	172 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	72 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_2_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_2_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_addr_2_ack_1, ack => testConfigure_CP_279_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	65 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	71 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_3_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_3_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_addr_3_ack_0, ack => testConfigure_CP_279_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	172 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	72 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_3_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_3_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_addr_3_ack_1, ack => testConfigure_CP_279_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	70 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_0/$exit
      -- CP-element group 81: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_store_0_ack_0, ack => testConfigure_CP_279_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_1/$exit
      -- CP-element group 82: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_1/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_store_1_ack_0, ack => testConfigure_CP_279_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	70 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_2/$exit
      -- CP-element group 83: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_2/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_store_2_ack_0, ack => testConfigure_CP_279_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	70 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_3/$exit
      -- CP-element group 84: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/word_3/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_store_3_ack_0, ack => testConfigure_CP_279_elements(84)); -- 
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	119 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(85) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(81) & testConfigure_CP_279_elements(82) & testConfigure_CP_279_elements(83) & testConfigure_CP_279_elements(84);
      gj_testConfigure_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	172 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	90 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_0/$exit
      -- CP-element group 86: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_store_0_ack_1, ack => testConfigure_CP_279_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	172 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_1/$exit
      -- CP-element group 87: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_1/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_store_1_ack_1, ack => testConfigure_CP_279_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	172 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_2/$exit
      -- CP-element group 88: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_2/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_store_2_ack_1, ack => testConfigure_CP_279_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	172 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_3/$exit
      -- CP-element group 89: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_3/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_184_store_3_ack_1, ack => testConfigure_CP_279_elements(89)); -- 
    -- CP-element group 90:  join  transition  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	86 
    -- CP-element group 90: 	87 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	120 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(90) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(86) & testConfigure_CP_279_elements(87) & testConfigure_CP_279_elements(88) & testConfigure_CP_279_elements(89);
      gj_testConfigure_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	67 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_update_start_
      -- CP-element group 91: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_Update/cr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:RPIPE_maxpool_input_pipe_188_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:RPIPE_maxpool_input_pipe_188_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_188_inst_ack_0, ack => testConfigure_CP_279_elements(91)); -- 
    cr_975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(91), ack => RPIPE_maxpool_input_pipe_188_inst_req_1); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_188_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_Sample/rr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:RPIPE_maxpool_input_pipe_188_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_192_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_188_inst_ack_1, ack => testConfigure_CP_279_elements(92)); -- 
    rr_984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(92), ack => type_cast_192_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_192_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_192_inst_ack_0, ack => testConfigure_CP_279_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	172 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_192_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_192_inst_ack_1, ack => testConfigure_CP_279_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: 	59 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/ptr_deref_195_Split/$entry
      -- CP-element group 95: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/ptr_deref_195_Split/$exit
      -- CP-element group 95: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/ptr_deref_195_Split/split_req
      -- CP-element group 95: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/ptr_deref_195_Split/split_ack
      -- CP-element group 95: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/word_access_start/$entry
      -- CP-element group 95: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/word_access_start/word_0/$entry
      -- CP-element group 95: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_195_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(95), ack => ptr_deref_195_store_0_req_0); -- 
    testConfigure_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(94) & testConfigure_CP_279_elements(59);
      gj_testConfigure_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/word_access_start/$exit
      -- CP-element group 96: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/word_access_start/word_0/$exit
      -- CP-element group 96: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_195_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_195_store_0_ack_0, ack => testConfigure_CP_279_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	172 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	120 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Update/word_access_complete/word_0/ca
      -- CP-element group 97: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Update/word_access_complete/word_0/$exit
      -- CP-element group 97: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Update/word_access_complete/$exit
      -- CP-element group 97: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_update_completed_
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_195_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_195_store_0_ack_1, ack => testConfigure_CP_279_elements(97)); -- 
    -- CP-element group 98:  join  fork  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	100 
    -- CP-element group 98: 	119 
    -- CP-element group 98: 	172 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	109 
    -- CP-element group 98: 	110 
    -- CP-element group 98: 	111 
    -- CP-element group 98: 	112 
    -- CP-element group 98:  members (11) 
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_3/rr
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_3/$entry
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_2/rr
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_2/$entry
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_1/rr
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_1/$entry
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_0/rr
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/$entry
      -- CP-element group 98: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_3_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(98), ack => ptr_deref_212_load_0_req_0); -- 
    rr_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(98), ack => ptr_deref_212_load_1_req_0); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(98), ack => ptr_deref_212_load_2_req_0); -- 
    rr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(98), ack => ptr_deref_212_load_3_req_0); -- 
    testConfigure_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(100) & testConfigure_CP_279_elements(119) & testConfigure_CP_279_elements(172);
      gj_testConfigure_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  join  transition  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	107 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	103 
    -- CP-element group 99: 	105 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	120 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_sample_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(99) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(107) & testConfigure_CP_279_elements(101) & testConfigure_CP_279_elements(103) & testConfigure_CP_279_elements(105);
      gj_testConfigure_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	108 
    -- CP-element group 100: 	102 
    -- CP-element group 100: 	104 
    -- CP-element group 100: 	106 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	98 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_address_calculated
      -- CP-element group 100: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_update_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(100) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(108) & testConfigure_CP_279_elements(102) & testConfigure_CP_279_elements(104) & testConfigure_CP_279_elements(106);
      gj_testConfigure_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	172 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	99 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_0_Sample/ra
      -- CP-element group 101: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_0_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_addr_0_ack_0, ack => testConfigure_CP_279_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	172 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	100 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_0_Update/ca
      -- CP-element group 102: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_0_Update/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_addr_0_ack_1, ack => testConfigure_CP_279_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	172 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	99 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_1_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_1_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(103) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_addr_1_ack_0, ack => testConfigure_CP_279_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	172 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	100 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_1_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_1_Update/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_addr_1_ack_1, ack => testConfigure_CP_279_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	172 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	99 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_2_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_2_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_addr_2_ack_0, ack => testConfigure_CP_279_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	172 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	100 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_2_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_2_Update/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_addr_2_ack_1, ack => testConfigure_CP_279_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	172 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	99 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_3_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_3_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_addr_3_ack_0, ack => testConfigure_CP_279_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	172 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	100 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_3_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_3_Update/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_addr_3_ack_1, ack => testConfigure_CP_279_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	98 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	113 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_0/ra
      -- CP-element group 109: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_0/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_load_0_ack_0, ack => testConfigure_CP_279_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	98 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_1/ra
      -- CP-element group 110: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_1/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_load_1_ack_0, ack => testConfigure_CP_279_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	98 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_2/ra
      -- CP-element group 111: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_2/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_load_2_ack_0, ack => testConfigure_CP_279_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	98 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_3/ra
      -- CP-element group 112: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/word_3/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_load_3_ack_0, ack => testConfigure_CP_279_elements(112)); -- 
    -- CP-element group 113:  join  transition  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	109 
    -- CP-element group 113: 	110 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/word_access_start/$exit
      -- CP-element group 113: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(113) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(109) & testConfigure_CP_279_elements(110) & testConfigure_CP_279_elements(111) & testConfigure_CP_279_elements(112);
      gj_testConfigure_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	172 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_0/$exit
      -- CP-element group 114: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_load_0_ack_1, ack => testConfigure_CP_279_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	172 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	118 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_1/ca
      -- CP-element group 115: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_1/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_load_1_ack_1, ack => testConfigure_CP_279_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	172 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_2/ca
      -- CP-element group 116: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_2/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_load_2_ack_1, ack => testConfigure_CP_279_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	172 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_3/ca
      -- CP-element group 117: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_3/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_212_load_3_ack_1, ack => testConfigure_CP_279_elements(117)); -- 
    -- CP-element group 118:  join  transition  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	115 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (7) 
      -- CP-element group 118: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/ptr_deref_212_Merge/$entry
      -- CP-element group 118: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/ptr_deref_212_Merge/merge_ack
      -- CP-element group 118: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/ptr_deref_212_Merge/merge_req
      -- CP-element group 118: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/ptr_deref_212_Merge/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(118) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(114) & testConfigure_CP_279_elements(115) & testConfigure_CP_279_elements(116) & testConfigure_CP_279_elements(117);
      gj_testConfigure_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  delay-element  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	85 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	98 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_ptr_deref_212_delay
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(119) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group testConfigure_CP_279_elements(119) is a control-delay.
    cp_element_119_delay: control_delay_element  generic map(name => " 119_delay", delay_value => 1)  port map(req => testConfigure_CP_279_elements(85), ack => testConfigure_CP_279_elements(119), clk => clk, reset =>reset);
    -- CP-element group 120:  branch  join  transition  place  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	56 
    -- CP-element group 120: 	60 
    -- CP-element group 120: 	62 
    -- CP-element group 120: 	99 
    -- CP-element group 120: 	71 
    -- CP-element group 120: 	97 
    -- CP-element group 120: 	90 
    -- CP-element group 120: 	55 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (10) 
      -- CP-element group 120: 	 branch_block_stmt_79/if_stmt_219_else_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_79/if_stmt_219_if_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_79/R_cmp_220_place
      -- CP-element group 120: 	 branch_block_stmt_79/if_stmt_219_eval_test/branch_req
      -- CP-element group 120: 	 branch_block_stmt_79/if_stmt_219_eval_test/$exit
      -- CP-element group 120: 	 branch_block_stmt_79/if_stmt_219_eval_test/$entry
      -- CP-element group 120: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/$exit
      -- CP-element group 120: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218__exit__
      -- CP-element group 120: 	 branch_block_stmt_79/if_stmt_219__entry__
      -- CP-element group 120: 	 branch_block_stmt_79/if_stmt_219_dead_link/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_219_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(120), ack => if_stmt_219_branch_req_0); -- 
    testConfigure_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(56) & testConfigure_CP_279_elements(60) & testConfigure_CP_279_elements(62) & testConfigure_CP_279_elements(99) & testConfigure_CP_279_elements(71) & testConfigure_CP_279_elements(97) & testConfigure_CP_279_elements(90) & testConfigure_CP_279_elements(55) & testConfigure_CP_279_elements(118);
      gj_testConfigure_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	168 
    -- CP-element group 121: 	169 
    -- CP-element group 121:  members (12) 
      -- CP-element group 121: 	 branch_block_stmt_79/if_stmt_219_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_79/if_stmt_219_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_79/forx_xbody_forx_xbody
      -- CP-element group 121: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/$entry
      -- CP-element group 121: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/$entry
      -- CP-element group 121: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/$entry
      -- CP-element group 121: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/SplitProtocol/$entry
      -- CP-element group 121: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/SplitProtocol/Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/SplitProtocol/Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/SplitProtocol/Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_219_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_150_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_150_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_219_branch_ack_1, ack => testConfigure_CP_279_elements(121)); -- 
    rr_1532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(121), ack => type_cast_150_inst_req_0); -- 
    cr_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(121), ack => type_cast_150_inst_req_1); -- 
    -- CP-element group 122:  fork  transition  place  input  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	163 
    -- CP-element group 122: 	164 
    -- CP-element group 122:  members (12) 
      -- CP-element group 122: 	 branch_block_stmt_79/if_stmt_219_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_79/if_stmt_219_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader
      -- CP-element group 122: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/$entry
      -- CP-element group 122: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/$entry
      -- CP-element group 122: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/$entry
      -- CP-element group 122: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/SplitProtocol/$entry
      -- CP-element group 122: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/SplitProtocol/Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/SplitProtocol/Sample/rr
      -- CP-element group 122: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/SplitProtocol/Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(122) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_219_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_129_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_129_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_219_branch_ack_0, ack => testConfigure_CP_279_elements(122)); -- 
    rr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(122), ack => type_cast_129_inst_req_0); -- 
    cr_1491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(122), ack => type_cast_129_inst_req_1); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	53 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_Sample/ra
      -- CP-element group 123: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_240_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_240_inst_ack_0, ack => testConfigure_CP_279_elements(123)); -- 
    -- CP-element group 124:  fork  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	53 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	173 
    -- CP-element group 124: 	174 
    -- CP-element group 124:  members (11) 
      -- CP-element group 124: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/$exit
      -- CP-element group 124: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254__exit__
      -- CP-element group 124: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18
      -- CP-element group 124: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_79/assign_stmt_231_to_assign_stmt_254/type_cast_240_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_257/$entry
      -- CP-element group 124: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_264/$entry
      -- CP-element group 124: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_240_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_240_inst_ack_1, ack => testConfigure_CP_279_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	186 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	152 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_276_index_1_scale_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_276_index_1_scale_ack_0, ack => testConfigure_CP_279_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	186 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (6) 
      -- CP-element group 126: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_update_complete
      -- CP-element group 126: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_final_index_sum_regn_Sample/req
      -- CP-element group 126: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_final_index_sum_regn_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scaled_1
      -- CP-element group 126: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_Update/ca
      -- CP-element group 126: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_Update/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_276_index_1_scale_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_276_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_276_index_1_scale_ack_1, ack => testConfigure_CP_279_elements(126)); -- 
    req_1233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(126), ack => array_obj_ref_276_index_offset_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	152 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_final_index_sum_regn_Sample/ack
      -- CP-element group 127: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_final_index_sum_regn_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_final_index_sum_regn_sample_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_276_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_276_index_offset_ack_0, ack => testConfigure_CP_279_elements(127)); -- 
    -- CP-element group 128:  transition  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	186 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (11) 
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_request/$entry
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_final_index_sum_regn_Update/ack
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_final_index_sum_regn_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_offset_calculated
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_request/req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_276_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_277_final_reg_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_276_index_offset_ack_1, ack => testConfigure_CP_279_elements(128)); -- 
    req_1248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(128), ack => addr_of_277_final_reg_req_0); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_request/ack
      -- CP-element group 129: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_request/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_277_final_reg_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_277_final_reg_ack_0, ack => testConfigure_CP_279_elements(129)); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	186 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	134 
    -- CP-element group 130: 	136 
    -- CP-element group 130: 	138 
    -- CP-element group 130: 	140 
    -- CP-element group 130:  members (23) 
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_sample_start
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_base_addr_resize/$exit
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_base_addr_resize/$entry
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_base_address_resized
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_root_address_calculated
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_base_plus_offset/sum_rename_ack
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_complete/ack
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_base_plus_offset/sum_rename_req
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_complete/$exit
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_1_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_0_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_base_address_calculated
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_0_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_1_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_base_plus_offset/$exit
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_base_plus_offset/$entry
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_3_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_3_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_base_addr_resize/base_resize_ack
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_2_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_2_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_base_addr_resize/base_resize_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_277_final_reg_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_3_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_277_final_reg_ack_1, ack => testConfigure_CP_279_elements(130)); -- 
    rr_1280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(130), ack => ptr_deref_281_addr_0_req_0); -- 
    rr_1290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(130), ack => ptr_deref_281_addr_1_req_0); -- 
    rr_1300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(130), ack => ptr_deref_281_addr_2_req_0); -- 
    rr_1310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(130), ack => ptr_deref_281_addr_3_req_0); -- 
    -- CP-element group 131:  join  fork  transition  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	142 
    -- CP-element group 131: 	143 
    -- CP-element group 131: 	144 
    -- CP-element group 131: 	145 
    -- CP-element group 131:  members (11) 
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_2/rr
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_2/$entry
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_1/rr
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_1/$entry
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_0/rr
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_0/$entry
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_3/rr
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/$entry
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_3/$entry
      -- CP-element group 131: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_sample_start_
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(131) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_3_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(131), ack => ptr_deref_281_load_0_req_0); -- 
    rr_1331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(131), ack => ptr_deref_281_load_1_req_0); -- 
    rr_1336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(131), ack => ptr_deref_281_load_2_req_0); -- 
    rr_1341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(131), ack => ptr_deref_281_load_3_req_0); -- 
    testConfigure_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(130) & testConfigure_CP_279_elements(133);
      gj_testConfigure_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: 	136 
    -- CP-element group 132: 	138 
    -- CP-element group 132: 	140 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	152 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_sample_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(132) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(134) & testConfigure_CP_279_elements(136) & testConfigure_CP_279_elements(138) & testConfigure_CP_279_elements(140);
      gj_testConfigure_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: 	137 
    -- CP-element group 133: 	139 
    -- CP-element group 133: 	141 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (2) 
      -- CP-element group 133: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_update_complete
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(133) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(135) & testConfigure_CP_279_elements(137) & testConfigure_CP_279_elements(139) & testConfigure_CP_279_elements(141);
      gj_testConfigure_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	130 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_0_Sample/ra
      -- CP-element group 134: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_0_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(134) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_addr_0_ack_0, ack => testConfigure_CP_279_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	186 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_0_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_0_Update/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(135) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_addr_0_ack_1, ack => testConfigure_CP_279_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	130 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	132 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_1_Sample/ra
      -- CP-element group 136: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_1_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(136) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_addr_1_ack_0, ack => testConfigure_CP_279_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	186 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	133 
    -- CP-element group 137:  members (2) 
      -- CP-element group 137: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_1_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_1_Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(137) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_addr_1_ack_1, ack => testConfigure_CP_279_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	130 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	132 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_2_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_2_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_addr_2_ack_0, ack => testConfigure_CP_279_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	186 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	133 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_2_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_2_Update/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(139) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_addr_2_ack_1, ack => testConfigure_CP_279_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	130 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	132 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_3_Sample/ra
      -- CP-element group 140: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_3_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_addr_3_ack_0, ack => testConfigure_CP_279_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	186 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	133 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_3_Update/ca
      -- CP-element group 141: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_3_Update/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(141) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_addr_3_ack_1, ack => testConfigure_CP_279_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	131 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	146 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_0/ra
      -- CP-element group 142: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_0/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(142) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_load_0_ack_0, ack => testConfigure_CP_279_elements(142)); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	131 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	146 
    -- CP-element group 143:  members (2) 
      -- CP-element group 143: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_1/ra
      -- CP-element group 143: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_1/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(143) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_load_1_ack_0, ack => testConfigure_CP_279_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	131 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_2/ra
      -- CP-element group 144: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_2/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(144) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_2_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_load_2_ack_0, ack => testConfigure_CP_279_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	131 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_3/ra
      -- CP-element group 145: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/word_3/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(145) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_3_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_load_3_ack_0, ack => testConfigure_CP_279_elements(145)); -- 
    -- CP-element group 146:  join  transition  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	142 
    -- CP-element group 146: 	143 
    -- CP-element group 146: 	144 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/word_access_start/$exit
      -- CP-element group 146: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_sample_completed_
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(146) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(142) & testConfigure_CP_279_elements(143) & testConfigure_CP_279_elements(144) & testConfigure_CP_279_elements(145);
      gj_testConfigure_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	186 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	151 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_0/ca
      -- CP-element group 147: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_0/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(147) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_load_0_ack_1, ack => testConfigure_CP_279_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	186 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	151 
    -- CP-element group 148:  members (2) 
      -- CP-element group 148: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_1/ca
      -- CP-element group 148: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_1/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(148) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_load_1_ack_1, ack => testConfigure_CP_279_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	186 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_2/$exit
      -- CP-element group 149: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_2/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(149) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_2_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_load_2_ack_1, ack => testConfigure_CP_279_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	186 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (2) 
      -- CP-element group 150: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_3/ca
      -- CP-element group 150: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_3/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(150) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_3_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_281_load_3_ack_1, ack => testConfigure_CP_279_elements(150)); -- 
    -- CP-element group 151:  join  transition  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	147 
    -- CP-element group 151: 	148 
    -- CP-element group 151: 	149 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (7) 
      -- CP-element group 151: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/$exit
      -- CP-element group 151: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/ptr_deref_281_Merge/merge_ack
      -- CP-element group 151: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/ptr_deref_281_Merge/$entry
      -- CP-element group 151: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/ptr_deref_281_Merge/$exit
      -- CP-element group 151: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/ptr_deref_281_Merge/merge_req
      -- CP-element group 151: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_update_completed_
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(151) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(147) & testConfigure_CP_279_elements(148) & testConfigure_CP_279_elements(149) & testConfigure_CP_279_elements(150);
      gj_testConfigure_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  branch  join  transition  place  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	125 
    -- CP-element group 152: 	127 
    -- CP-element group 152: 	132 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (10) 
      -- CP-element group 152: 	 branch_block_stmt_79/if_stmt_299_eval_test/branch_req
      -- CP-element group 152: 	 branch_block_stmt_79/R_exitcond_300_place
      -- CP-element group 152: 	 branch_block_stmt_79/if_stmt_299_dead_link/$entry
      -- CP-element group 152: 	 branch_block_stmt_79/if_stmt_299_eval_test/$entry
      -- CP-element group 152: 	 branch_block_stmt_79/if_stmt_299_eval_test/$exit
      -- CP-element group 152: 	 branch_block_stmt_79/if_stmt_299_if_link/$entry
      -- CP-element group 152: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298__exit__
      -- CP-element group 152: 	 branch_block_stmt_79/if_stmt_299__entry__
      -- CP-element group 152: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/$exit
      -- CP-element group 152: 	 branch_block_stmt_79/if_stmt_299_else_link/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(152) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_299_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(152), ack => if_stmt_299_branch_req_0); -- 
    testConfigure_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(125) & testConfigure_CP_279_elements(127) & testConfigure_CP_279_elements(132) & testConfigure_CP_279_elements(151);
      gj_testConfigure_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  place  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	187 
    -- CP-element group 153: 	188 
    -- CP-element group 153: 	190 
    -- CP-element group 153: 	191 
    -- CP-element group 153: 	193 
    -- CP-element group 153: 	194 
    -- CP-element group 153:  members (28) 
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27
      -- CP-element group 153: 	 branch_block_stmt_79/if_stmt_299_if_link/$exit
      -- CP-element group 153: 	 branch_block_stmt_79/if_stmt_299_if_link/if_choice_transition
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/SplitProtocol/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/SplitProtocol/Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/SplitProtocol/Sample/rr
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/SplitProtocol/Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/SplitProtocol/Update/cr
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/rr
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/cr
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/SplitProtocol/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/SplitProtocol/Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/SplitProtocol/Sample/rr
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/SplitProtocol/Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(153) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_299_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_313_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_313_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_309_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_309_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_317_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_317_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_299_branch_ack_1, ack => testConfigure_CP_279_elements(153)); -- 
    rr_1653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(153), ack => type_cast_313_inst_req_0); -- 
    cr_1658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(153), ack => type_cast_313_inst_req_1); -- 
    rr_1676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(153), ack => type_cast_309_inst_req_0); -- 
    cr_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(153), ack => type_cast_309_inst_req_1); -- 
    rr_1699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(153), ack => type_cast_317_inst_req_0); -- 
    cr_1704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(153), ack => type_cast_317_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  place  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	176 
    -- CP-element group 154: 	177 
    -- CP-element group 154: 	179 
    -- CP-element group 154: 	180 
    -- CP-element group 154:  members (20) 
      -- CP-element group 154: 	 branch_block_stmt_79/if_stmt_299_else_link/else_choice_transition
      -- CP-element group 154: 	 branch_block_stmt_79/if_stmt_299_else_link/$exit
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/cr
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/SplitProtocol/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/SplitProtocol/Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/SplitProtocol/Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/SplitProtocol/Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(154) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_299_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_263_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_263_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_270_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_270_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_299_branch_ack_0, ack => testConfigure_CP_279_elements(154)); -- 
    rr_1594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(154), ack => type_cast_263_inst_req_0); -- 
    cr_1599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(154), ack => type_cast_263_inst_req_1); -- 
    rr_1617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(154), ack => type_cast_270_inst_req_0); -- 
    cr_1622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(154), ack => type_cast_270_inst_req_1); -- 
    -- CP-element group 155:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	1 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: 	158 
    -- CP-element group 155:  members (18) 
      -- CP-element group 155: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/$entry
      -- CP-element group 155: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_update_start_
      -- CP-element group 155: 	 branch_block_stmt_79/if_stmt_325_if_link/if_choice_transition
      -- CP-element group 155: 	 branch_block_stmt_79/if_stmt_325_if_link/$exit
      -- CP-element group 155: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_Update/cr
      -- CP-element group 155: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_79/forx_xend27_bbx_xnph
      -- CP-element group 155: 	 branch_block_stmt_79/merge_stmt_331__exit__
      -- CP-element group 155: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361__entry__
      -- CP-element group 155: 	 branch_block_stmt_79/forx_xend27_bbx_xnph_PhiReq/$entry
      -- CP-element group 155: 	 branch_block_stmt_79/forx_xend27_bbx_xnph_PhiReq/$exit
      -- CP-element group 155: 	 branch_block_stmt_79/merge_stmt_331_PhiReqMerge
      -- CP-element group 155: 	 branch_block_stmt_79/merge_stmt_331_PhiAck/$entry
      -- CP-element group 155: 	 branch_block_stmt_79/merge_stmt_331_PhiAck/$exit
      -- CP-element group 155: 	 branch_block_stmt_79/merge_stmt_331_PhiAck/dummy
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(155) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_325_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_341_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_341_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_325_branch_ack_1, ack => testConfigure_CP_279_elements(155)); -- 
    rr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(155), ack => type_cast_341_inst_req_0); -- 
    cr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(155), ack => type_cast_341_inst_req_1); -- 
    -- CP-element group 156:  transition  place  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	1 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	207 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_79/if_stmt_325_else_link/$exit
      -- CP-element group 156: 	 branch_block_stmt_79/if_stmt_325_else_link/else_choice_transition
      -- CP-element group 156: 	 branch_block_stmt_79/forx_xend27_forx_xend42
      -- CP-element group 156: 	 branch_block_stmt_79/forx_xend27_forx_xend42_PhiReq/$entry
      -- CP-element group 156: 	 branch_block_stmt_79/forx_xend27_forx_xend42_PhiReq/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_325_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_325_branch_ack_0, ack => testConfigure_CP_279_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_Sample/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_341_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_341_inst_ack_0, ack => testConfigure_CP_279_elements(157)); -- 
    -- CP-element group 158:  transition  place  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	155 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	201 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/$exit
      -- CP-element group 158: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361/type_cast_341_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_79/assign_stmt_336_to_assign_stmt_361__exit__
      -- CP-element group 158: 	 branch_block_stmt_79/bbx_xnph_forx_xbody36
      -- CP-element group 158: 	 branch_block_stmt_79/bbx_xnph_forx_xbody36_PhiReq/$entry
      -- CP-element group 158: 	 branch_block_stmt_79/bbx_xnph_forx_xbody36_PhiReq/phi_stmt_364/$entry
      -- CP-element group 158: 	 branch_block_stmt_79/bbx_xnph_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(158) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_341_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_341_inst_ack_1, ack => testConfigure_CP_279_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	206 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_Sample/cra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:call_stmt_373_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_373_call_ack_0, ack => testConfigure_CP_279_elements(159)); -- 
    -- CP-element group 160:  branch  transition  place  input  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	206 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (13) 
      -- CP-element group 160: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/$exit
      -- CP-element group 160: 	 branch_block_stmt_79/if_stmt_385_dead_link/$entry
      -- CP-element group 160: 	 branch_block_stmt_79/if_stmt_385_else_link/$entry
      -- CP-element group 160: 	 branch_block_stmt_79/R_exitcond7_386_place
      -- CP-element group 160: 	 branch_block_stmt_79/if_stmt_385_if_link/$entry
      -- CP-element group 160: 	 branch_block_stmt_79/if_stmt_385_eval_test/$entry
      -- CP-element group 160: 	 branch_block_stmt_79/if_stmt_385_eval_test/$exit
      -- CP-element group 160: 	 branch_block_stmt_79/if_stmt_385_eval_test/branch_req
      -- CP-element group 160: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_Update/cca
      -- CP-element group 160: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384__exit__
      -- CP-element group 160: 	 branch_block_stmt_79/if_stmt_385__entry__
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(160) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:call_stmt_373_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_385_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_1448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_373_call_ack_1, ack => testConfigure_CP_279_elements(160)); -- 
    branch_req_1456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(160), ack => if_stmt_385_branch_req_0); -- 
    -- CP-element group 161:  merge  transition  place  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	207 
    -- CP-element group 161:  members (13) 
      -- CP-element group 161: 	 branch_block_stmt_79/if_stmt_385_if_link/if_choice_transition
      -- CP-element group 161: 	 branch_block_stmt_79/if_stmt_385_if_link/$exit
      -- CP-element group 161: 	 branch_block_stmt_79/forx_xbody36_forx_xend42x_xloopexit
      -- CP-element group 161: 	 branch_block_stmt_79/merge_stmt_391__exit__
      -- CP-element group 161: 	 branch_block_stmt_79/forx_xend42x_xloopexit_forx_xend42
      -- CP-element group 161: 	 branch_block_stmt_79/forx_xbody36_forx_xend42x_xloopexit_PhiReq/$entry
      -- CP-element group 161: 	 branch_block_stmt_79/forx_xbody36_forx_xend42x_xloopexit_PhiReq/$exit
      -- CP-element group 161: 	 branch_block_stmt_79/merge_stmt_391_PhiReqMerge
      -- CP-element group 161: 	 branch_block_stmt_79/merge_stmt_391_PhiAck/$entry
      -- CP-element group 161: 	 branch_block_stmt_79/merge_stmt_391_PhiAck/$exit
      -- CP-element group 161: 	 branch_block_stmt_79/merge_stmt_391_PhiAck/dummy
      -- CP-element group 161: 	 branch_block_stmt_79/forx_xend42x_xloopexit_forx_xend42_PhiReq/$entry
      -- CP-element group 161: 	 branch_block_stmt_79/forx_xend42x_xloopexit_forx_xend42_PhiReq/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(161) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_385_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_385_branch_ack_1, ack => testConfigure_CP_279_elements(161)); -- 
    -- CP-element group 162:  fork  transition  place  input  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	202 
    -- CP-element group 162: 	203 
    -- CP-element group 162:  members (12) 
      -- CP-element group 162: 	 branch_block_stmt_79/if_stmt_385_else_link/$exit
      -- CP-element group 162: 	 branch_block_stmt_79/if_stmt_385_else_link/else_choice_transition
      -- CP-element group 162: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36
      -- CP-element group 162: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/$entry
      -- CP-element group 162: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/$entry
      -- CP-element group 162: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/$entry
      -- CP-element group 162: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/$entry
      -- CP-element group 162: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/SplitProtocol/$entry
      -- CP-element group 162: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/SplitProtocol/Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/SplitProtocol/Sample/rr
      -- CP-element group 162: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/SplitProtocol/Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/SplitProtocol/Update/cr
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_385_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_370_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_370_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_385_branch_ack_0, ack => testConfigure_CP_279_elements(162)); -- 
    rr_1755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(162), ack => type_cast_370_inst_req_0); -- 
    cr_1760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(162), ack => type_cast_370_inst_req_1); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	122 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/SplitProtocol/Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_129_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_129_inst_ack_0, ack => testConfigure_CP_279_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	122 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/SplitProtocol/Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(164) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_129_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_129_inst_ack_1, ack => testConfigure_CP_279_elements(164)); -- 
    -- CP-element group 165:  join  transition  place  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (8) 
      -- CP-element group 165: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/$exit
      -- CP-element group 165: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/$exit
      -- CP-element group 165: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/$exit
      -- CP-element group 165: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_sources/type_cast_129/SplitProtocol/$exit
      -- CP-element group 165: 	 branch_block_stmt_79/forx_xbody_forx_xcond13x_xpreheader_PhiReq/phi_stmt_126/phi_stmt_126_req
      -- CP-element group 165: 	 branch_block_stmt_79/merge_stmt_125_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_79/merge_stmt_125_PhiAck/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_126_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_126_req_1493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_126_req_1493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(165), ack => phi_stmt_126_req_0); -- 
    testConfigure_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(163) & testConfigure_CP_279_elements(164);
      gj_testConfigure_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  branch  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	52 
    -- CP-element group 166: 	53 
    -- CP-element group 166:  members (15) 
      -- CP-element group 166: 	 branch_block_stmt_79/assign_stmt_136/$entry
      -- CP-element group 166: 	 branch_block_stmt_79/assign_stmt_136/$exit
      -- CP-element group 166: 	 branch_block_stmt_79/if_stmt_137_dead_link/$entry
      -- CP-element group 166: 	 branch_block_stmt_79/if_stmt_137_eval_test/$entry
      -- CP-element group 166: 	 branch_block_stmt_79/if_stmt_137_eval_test/$exit
      -- CP-element group 166: 	 branch_block_stmt_79/if_stmt_137_eval_test/branch_req
      -- CP-element group 166: 	 branch_block_stmt_79/R_cmp1648_138_place
      -- CP-element group 166: 	 branch_block_stmt_79/if_stmt_137_if_link/$entry
      -- CP-element group 166: 	 branch_block_stmt_79/if_stmt_137_else_link/$entry
      -- CP-element group 166: 	 branch_block_stmt_79/merge_stmt_125__exit__
      -- CP-element group 166: 	 branch_block_stmt_79/assign_stmt_136__entry__
      -- CP-element group 166: 	 branch_block_stmt_79/assign_stmt_136__exit__
      -- CP-element group 166: 	 branch_block_stmt_79/if_stmt_137__entry__
      -- CP-element group 166: 	 branch_block_stmt_79/merge_stmt_125_PhiAck/$exit
      -- CP-element group 166: 	 branch_block_stmt_79/merge_stmt_125_PhiAck/phi_stmt_126_ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(166) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_126_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:if_stmt_137_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_126_ack_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_126_ack_0, ack => testConfigure_CP_279_elements(166)); -- 
    branch_req_686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(166), ack => if_stmt_137_branch_req_0); -- 
    -- CP-element group 167:  transition  output  delay-element  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	51 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	171 
    -- CP-element group 167:  members (5) 
      -- CP-element group 167: 	 branch_block_stmt_79/bbx_xnph55_forx_xbody_PhiReq/$exit
      -- CP-element group 167: 	 branch_block_stmt_79/bbx_xnph55_forx_xbody_PhiReq/phi_stmt_144/$exit
      -- CP-element group 167: 	 branch_block_stmt_79/bbx_xnph55_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/$exit
      -- CP-element group 167: 	 branch_block_stmt_79/bbx_xnph55_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_148_konst_delay_trans
      -- CP-element group 167: 	 branch_block_stmt_79/bbx_xnph55_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_144_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_144_req_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_144_req_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(167), ack => phi_stmt_144_req_0); -- 
    -- Element group testConfigure_CP_279_elements(167) is a control-delay.
    cp_element_167_delay: control_delay_element  generic map(name => " 167_delay", delay_value => 1)  port map(req => testConfigure_CP_279_elements(51), ack => testConfigure_CP_279_elements(167), clk => clk, reset =>reset);
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (2) 
      -- CP-element group 168: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/SplitProtocol/Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(168)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(168)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(168) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_150_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_150_inst_ack_0, ack => testConfigure_CP_279_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	121 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (2) 
      -- CP-element group 169: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/SplitProtocol/Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(169)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(169)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(169) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_150_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_150_inst_ack_1, ack => testConfigure_CP_279_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (6) 
      -- CP-element group 170: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 170: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/$exit
      -- CP-element group 170: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/$exit
      -- CP-element group 170: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/$exit
      -- CP-element group 170: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_150/SplitProtocol/$exit
      -- CP-element group 170: 	 branch_block_stmt_79/forx_xbody_forx_xbody_PhiReq/phi_stmt_144/phi_stmt_144_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(170)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(170)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(170) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_144_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_144_req_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_144_req_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(170), ack => phi_stmt_144_req_1); -- 
    testConfigure_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(168) & testConfigure_CP_279_elements(169);
      gj_testConfigure_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  merge  transition  place  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	167 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (2) 
      -- CP-element group 171: 	 branch_block_stmt_79/merge_stmt_143_PhiReqMerge
      -- CP-element group 171: 	 branch_block_stmt_79/merge_stmt_143_PhiAck/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(171)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(171)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(171) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_CP_279_elements(171) <= OrReduce(testConfigure_CP_279_elements(167) & testConfigure_CP_279_elements(170));
    -- CP-element group 172:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	56 
    -- CP-element group 172: 	57 
    -- CP-element group 172: 	94 
    -- CP-element group 172: 	59 
    -- CP-element group 172: 	60 
    -- CP-element group 172: 	61 
    -- CP-element group 172: 	63 
    -- CP-element group 172: 	107 
    -- CP-element group 172: 	108 
    -- CP-element group 172: 	65 
    -- CP-element group 172: 	101 
    -- CP-element group 172: 	66 
    -- CP-element group 172: 	69 
    -- CP-element group 172: 	74 
    -- CP-element group 172: 	76 
    -- CP-element group 172: 	97 
    -- CP-element group 172: 	98 
    -- CP-element group 172: 	78 
    -- CP-element group 172: 	80 
    -- CP-element group 172: 	86 
    -- CP-element group 172: 	87 
    -- CP-element group 172: 	88 
    -- CP-element group 172: 	102 
    -- CP-element group 172: 	103 
    -- CP-element group 172: 	104 
    -- CP-element group 172: 	105 
    -- CP-element group 172: 	106 
    -- CP-element group 172: 	89 
    -- CP-element group 172: 	54 
    -- CP-element group 172: 	55 
    -- CP-element group 172: 	114 
    -- CP-element group 172: 	115 
    -- CP-element group 172: 	116 
    -- CP-element group 172: 	117 
    -- CP-element group 172:  members (122) 
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_3_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_0/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_sample_start
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_3_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_3_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_3_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_update_start
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_update_start_
      -- CP-element group 172: 	 branch_block_stmt_79/merge_stmt_143__exit__
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218__entry__
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_2_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_2_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_update_start_
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_2_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_2_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_1_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_1_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_1_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_1_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Update/word_access_complete/word_0/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_0_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_0_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Update/word_access_complete/word_0/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_3/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_0_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_3/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_2/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_2/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_Update/word_access_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_word_addrgen_0_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_1/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_1/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_212_Update/word_access_complete/word_0/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_160_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_update_start_
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_resized_1
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_scaled_1
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_computed_1
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_resize_1/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_resize_1/$exit
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_resize_1/index_resize_req
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_resize_1/index_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_scale_1/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_scale_1/$exit
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_scale_1/scale_rename_req
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_index_scale_1/scale_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_final_index_sum_regn_update_start
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_final_index_sum_regn_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_final_index_sum_regn_Sample/req
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_final_index_sum_regn_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_166_final_index_sum_regn_Update/req
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_167_complete/req
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_update_start_
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_resized_1
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_computed_1
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_resize_1/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_resize_1/$exit
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_resize_1/index_resize_req
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_resize_1/index_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_sample_start
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_update_start
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_index_scale_1_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_final_index_sum_regn_update_start
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_final_index_sum_regn_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/array_obj_ref_173_final_index_sum_regn_Update/req
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/addr_of_174_complete/req
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/RPIPE_maxpool_input_pipe_177_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_update_start_
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_181_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_update_start_
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_update_start
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_0_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_0_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_1_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_1_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_2_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_2_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_3_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_word_addrgen_3_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_0/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_0/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_1/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_1/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_2/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_2/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_3/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_184_Update/word_access_complete/word_3/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_update_start_
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/type_cast_192_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_79/assign_stmt_157_to_assign_stmt_218/ptr_deref_195_update_start_
      -- CP-element group 172: 	 branch_block_stmt_79/merge_stmt_143_PhiAck/$exit
      -- CP-element group 172: 	 branch_block_stmt_79/merge_stmt_143_PhiAck/phi_stmt_144_ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(172)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(172)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(172) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_144_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_3_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_2_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_1_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_195_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_addr_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_212_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_160_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_160_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_166_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_166_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_167_final_reg_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_173_index_1_scale_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_173_index_1_scale_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_173_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_174_final_reg_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:RPIPE_maxpool_input_pipe_177_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_181_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_addr_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_184_store_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_192_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_144_ack_1544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_144_ack_0, ack => testConfigure_CP_279_elements(172)); -- 
    cr_1101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_addr_3_req_1); -- 
    rr_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_addr_3_req_0); -- 
    cr_1091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_addr_2_req_1); -- 
    rr_1086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_addr_2_req_0); -- 
    cr_1081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_addr_1_req_1); -- 
    rr_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_addr_1_req_0); -- 
    cr_1039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_195_store_0_req_1); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_addr_0_req_1); -- 
    cr_1153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_load_3_req_1); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_addr_0_req_0); -- 
    cr_1148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_load_2_req_1); -- 
    cr_1143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_load_1_req_1); -- 
    cr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_212_load_0_req_1); -- 
    rr_708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => type_cast_160_inst_req_0); -- 
    cr_713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => type_cast_160_inst_req_1); -- 
    req_739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => array_obj_ref_166_index_offset_req_0); -- 
    req_744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => array_obj_ref_166_index_offset_req_1); -- 
    req_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => addr_of_167_final_reg_req_1); -- 
    rr_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => array_obj_ref_173_index_1_scale_req_0); -- 
    cr_787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => array_obj_ref_173_index_1_scale_req_1); -- 
    req_799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => array_obj_ref_173_index_offset_req_1); -- 
    req_814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => addr_of_174_final_reg_req_1); -- 
    rr_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => RPIPE_maxpool_input_pipe_177_inst_req_0); -- 
    cr_842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => type_cast_181_inst_req_1); -- 
    cr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_184_addr_0_req_1); -- 
    cr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_184_addr_1_req_1); -- 
    cr_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_184_addr_2_req_1); -- 
    cr_904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_184_addr_3_req_1); -- 
    cr_946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_184_store_0_req_1); -- 
    cr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_184_store_1_req_1); -- 
    cr_956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_184_store_2_req_1); -- 
    cr_961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => ptr_deref_184_store_3_req_1); -- 
    cr_989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(172), ack => type_cast_192_inst_req_1); -- 
    -- CP-element group 173:  transition  output  delay-element  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	124 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (4) 
      -- CP-element group 173: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_257/$exit
      -- CP-element group 173: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/$exit
      -- CP-element group 173: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_261_konst_delay_trans
      -- CP-element group 173: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(173)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(173)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(173) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_257_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_257_req_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_257_req_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(173), ack => phi_stmt_257_req_0); -- 
    -- Element group testConfigure_CP_279_elements(173) is a control-delay.
    cp_element_173_delay: control_delay_element  generic map(name => " 173_delay", delay_value => 1)  port map(req => testConfigure_CP_279_elements(124), ack => testConfigure_CP_279_elements(173), clk => clk, reset =>reset);
    -- CP-element group 174:  transition  output  delay-element  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	124 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (4) 
      -- CP-element group 174: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_264/$exit
      -- CP-element group 174: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/$exit
      -- CP-element group 174: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_268_konst_delay_trans
      -- CP-element group 174: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(174)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(174)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(174) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_264_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_264_req_1575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_264_req_1575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(174), ack => phi_stmt_264_req_0); -- 
    -- Element group testConfigure_CP_279_elements(174) is a control-delay.
    cp_element_174_delay: control_delay_element  generic map(name => " 174_delay", delay_value => 1)  port map(req => testConfigure_CP_279_elements(124), ack => testConfigure_CP_279_elements(174), clk => clk, reset =>reset);
    -- CP-element group 175:  join  transition  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	183 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 branch_block_stmt_79/bbx_xnph51_forx_xbody18_PhiReq/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(175)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(175)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(175) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(173) & testConfigure_CP_279_elements(174);
      gj_testConfigure_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	154 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (2) 
      -- CP-element group 176: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(176)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(176)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(176) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_263_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_0, ack => testConfigure_CP_279_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	154 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (2) 
      -- CP-element group 177: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(177)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(177)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(177) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_263_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_1, ack => testConfigure_CP_279_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	182 
    -- CP-element group 178:  members (5) 
      -- CP-element group 178: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/$exit
      -- CP-element group 178: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/$exit
      -- CP-element group 178: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/$exit
      -- CP-element group 178: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/$exit
      -- CP-element group 178: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_257/phi_stmt_257_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(178)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(178)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(178) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_257_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_257_req_1601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_257_req_1601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(178), ack => phi_stmt_257_req_1); -- 
    testConfigure_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(176) & testConfigure_CP_279_elements(177);
      gj_testConfigure_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	154 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (2) 
      -- CP-element group 179: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/SplitProtocol/Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(179)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(179)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(179) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_270_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_270_inst_ack_0, ack => testConfigure_CP_279_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	154 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/SplitProtocol/Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(180)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(180)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(180) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_270_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_270_inst_ack_1, ack => testConfigure_CP_279_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/$exit
      -- CP-element group 181: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/$exit
      -- CP-element group 181: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/$exit
      -- CP-element group 181: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_270/SplitProtocol/$exit
      -- CP-element group 181: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/phi_stmt_264/phi_stmt_264_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(181)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(181)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(181) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_264_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_264_req_1624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_264_req_1624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(181), ack => phi_stmt_264_req_1); -- 
    testConfigure_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(179) & testConfigure_CP_279_elements(180);
      gj_testConfigure_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  join  transition  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	178 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_79/forx_xbody18_forx_xbody18_PhiReq/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(182)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(182)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(182) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(178) & testConfigure_CP_279_elements(181);
      gj_testConfigure_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  merge  fork  transition  place  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	175 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_79/merge_stmt_256_PhiReqMerge
      -- CP-element group 183: 	 branch_block_stmt_79/merge_stmt_256_PhiAck/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(183)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(183)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(183) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_CP_279_elements(183) <= OrReduce(testConfigure_CP_279_elements(175) & testConfigure_CP_279_elements(182));
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_79/merge_stmt_256_PhiAck/phi_stmt_257_ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(184)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(184)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(184) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_257_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_257_ack_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_257_ack_0, ack => testConfigure_CP_279_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_79/merge_stmt_256_PhiAck/phi_stmt_264_ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(185)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(185)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(185) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_264_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_264_ack_1630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_264_ack_0, ack => testConfigure_CP_279_elements(185)); -- 
    -- CP-element group 186:  join  fork  transition  place  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	125 
    -- CP-element group 186: 	126 
    -- CP-element group 186: 	128 
    -- CP-element group 186: 	130 
    -- CP-element group 186: 	135 
    -- CP-element group 186: 	137 
    -- CP-element group 186: 	139 
    -- CP-element group 186: 	141 
    -- CP-element group 186: 	147 
    -- CP-element group 186: 	148 
    -- CP-element group 186: 	149 
    -- CP-element group 186: 	150 
    -- CP-element group 186:  members (42) 
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_update_start
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_1_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_0_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_0/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_1_Update/cr
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_update_start
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_resize_1/index_resize_ack
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_sample_start
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_complete/req
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_final_index_sum_regn_Update/req
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_final_index_sum_regn_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_2/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_1/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_0_Update/cr
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_resize_1/index_resize_req
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_resize_1/$exit
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_resize_1/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_3/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_0/cr
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_final_index_sum_regn_update_start
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_1/cr
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_2/cr
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_complete/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_Update/word_access_complete/word_3/cr
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_computed_1
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_update_start_
      -- CP-element group 186: 	 branch_block_stmt_79/merge_stmt_256__exit__
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298__entry__
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_resized_1
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_3_Update/cr
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/addr_of_277_update_start_
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_3_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_Update/cr
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/array_obj_ref_276_index_scale_1_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_2_Update/cr
      -- CP-element group 186: 	 branch_block_stmt_79/assign_stmt_278_to_assign_stmt_298/ptr_deref_281_word_addrgen_2_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_79/merge_stmt_256_PhiAck/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(186)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(186)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(186) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:addr_of_277_final_reg_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_276_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_1_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_276_index_1_scale_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_2_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_load_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_3_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:array_obj_ref_276_index_1_scale_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:ptr_deref_281_addr_2_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => ptr_deref_281_addr_1_req_1); -- 
    req_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => addr_of_277_final_reg_req_1); -- 
    req_1238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => array_obj_ref_276_index_offset_req_1); -- 
    cr_1285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => ptr_deref_281_addr_0_req_1); -- 
    cr_1352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => ptr_deref_281_load_0_req_1); -- 
    cr_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => ptr_deref_281_load_1_req_1); -- 
    rr_1221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => array_obj_ref_276_index_1_scale_req_0); -- 
    cr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => ptr_deref_281_load_2_req_1); -- 
    cr_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => ptr_deref_281_load_3_req_1); -- 
    cr_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => ptr_deref_281_addr_3_req_1); -- 
    cr_1226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => array_obj_ref_276_index_1_scale_req_1); -- 
    cr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(186), ack => ptr_deref_281_addr_2_req_1); -- 
    testConfigure_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(184) & testConfigure_CP_279_elements(185);
      gj_testConfigure_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	153 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (2) 
      -- CP-element group 187: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/SplitProtocol/Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(187)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(187)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(187) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_313_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_313_inst_ack_0, ack => testConfigure_CP_279_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	153 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (2) 
      -- CP-element group 188: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/SplitProtocol/Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(188)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(188)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(188) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_313_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_313_inst_ack_1, ack => testConfigure_CP_279_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	196 
    -- CP-element group 189:  members (5) 
      -- CP-element group 189: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/$exit
      -- CP-element group 189: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/$exit
      -- CP-element group 189: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/$exit
      -- CP-element group 189: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_sources/type_cast_313/SplitProtocol/$exit
      -- CP-element group 189: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_310/phi_stmt_310_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(189)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(189)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(189) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_310_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_310_req_1660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_310_req_1660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(189), ack => phi_stmt_310_req_0); -- 
    testConfigure_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(187) & testConfigure_CP_279_elements(188);
      gj_testConfigure_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	153 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (2) 
      -- CP-element group 190: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(190)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(190)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(190) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_309_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_309_inst_ack_0, ack => testConfigure_CP_279_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	153 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (2) 
      -- CP-element group 191: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(191)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(191)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(191) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_309_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_309_inst_ack_1, ack => testConfigure_CP_279_elements(191)); -- 
    -- CP-element group 192:  join  transition  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	196 
    -- CP-element group 192:  members (5) 
      -- CP-element group 192: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/$exit
      -- CP-element group 192: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/$exit
      -- CP-element group 192: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/$exit
      -- CP-element group 192: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/$exit
      -- CP-element group 192: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_306/phi_stmt_306_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(192)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(192)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(192) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_306_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_306_req_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_306_req_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(192), ack => phi_stmt_306_req_0); -- 
    testConfigure_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(190) & testConfigure_CP_279_elements(191);
      gj_testConfigure_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	153 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (2) 
      -- CP-element group 193: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/SplitProtocol/Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(193)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(193)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(193) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_317_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_317_inst_ack_0, ack => testConfigure_CP_279_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	153 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (2) 
      -- CP-element group 194: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/SplitProtocol/Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(194)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(194)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(194) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_317_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_317_inst_ack_1, ack => testConfigure_CP_279_elements(194)); -- 
    -- CP-element group 195:  join  transition  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (5) 
      -- CP-element group 195: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/$exit
      -- CP-element group 195: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/$exit
      -- CP-element group 195: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/$exit
      -- CP-element group 195: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_sources/type_cast_317/SplitProtocol/$exit
      -- CP-element group 195: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/phi_stmt_314/phi_stmt_314_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(195)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(195)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(195) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_314_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_314_req_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_314_req_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(195), ack => phi_stmt_314_req_0); -- 
    testConfigure_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(193) & testConfigure_CP_279_elements(194);
      gj_testConfigure_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  join  fork  transition  place  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	189 
    -- CP-element group 196: 	192 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	198 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_79/forx_xbody18_forx_xend27_PhiReq/$exit
      -- CP-element group 196: 	 branch_block_stmt_79/merge_stmt_305_PhiReqMerge
      -- CP-element group 196: 	 branch_block_stmt_79/merge_stmt_305_PhiAck/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(196)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(196)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(196) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(189) & testConfigure_CP_279_elements(192) & testConfigure_CP_279_elements(195);
      gj_testConfigure_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	200 
    -- CP-element group 197:  members (1) 
      -- CP-element group 197: 	 branch_block_stmt_79/merge_stmt_305_PhiAck/phi_stmt_306_ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(197)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(197)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(197) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_306_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_306_ack_1711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_306_ack_0, ack => testConfigure_CP_279_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_79/merge_stmt_305_PhiAck/phi_stmt_310_ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(198)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(198)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(198) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_310_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_310_ack_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_310_ack_0, ack => testConfigure_CP_279_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (1) 
      -- CP-element group 199: 	 branch_block_stmt_79/merge_stmt_305_PhiAck/phi_stmt_314_ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(199)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(199)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(199) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_314_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_314_ack_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_314_ack_0, ack => testConfigure_CP_279_elements(199)); -- 
    -- CP-element group 200:  join  transition  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	197 
    -- CP-element group 200: 	198 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	1 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_79/merge_stmt_305_PhiAck/$exit
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(200)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(200)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(200) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(197) & testConfigure_CP_279_elements(198) & testConfigure_CP_279_elements(199);
      gj_testConfigure_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  transition  output  delay-element  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	158 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	205 
    -- CP-element group 201:  members (5) 
      -- CP-element group 201: 	 branch_block_stmt_79/bbx_xnph_forx_xbody36_PhiReq/$exit
      -- CP-element group 201: 	 branch_block_stmt_79/bbx_xnph_forx_xbody36_PhiReq/phi_stmt_364/$exit
      -- CP-element group 201: 	 branch_block_stmt_79/bbx_xnph_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/$exit
      -- CP-element group 201: 	 branch_block_stmt_79/bbx_xnph_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_368_konst_delay_trans
      -- CP-element group 201: 	 branch_block_stmt_79/bbx_xnph_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(201)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(201)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(201) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_364_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_364_req_1736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_364_req_1736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(201), ack => phi_stmt_364_req_0); -- 
    -- Element group testConfigure_CP_279_elements(201) is a control-delay.
    cp_element_201_delay: control_delay_element  generic map(name => " 201_delay", delay_value => 1)  port map(req => testConfigure_CP_279_elements(158), ack => testConfigure_CP_279_elements(201), clk => clk, reset =>reset);
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	162 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (2) 
      -- CP-element group 202: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/SplitProtocol/Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/SplitProtocol/Sample/ra
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(202)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(202)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(202) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_370_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_0, ack => testConfigure_CP_279_elements(202)); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	162 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (2) 
      -- CP-element group 203: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/SplitProtocol/Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/SplitProtocol/Update/ca
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(203)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(203)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(203) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:type_cast_370_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_1, ack => testConfigure_CP_279_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/$exit
      -- CP-element group 204: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/$exit
      -- CP-element group 204: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/$exit
      -- CP-element group 204: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/$exit
      -- CP-element group 204: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_sources/type_cast_370/SplitProtocol/$exit
      -- CP-element group 204: 	 branch_block_stmt_79/forx_xbody36_forx_xbody36_PhiReq/phi_stmt_364/phi_stmt_364_req
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(204)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(204)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(204) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_364_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_364_req_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_364_req_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(204), ack => phi_stmt_364_req_1); -- 
    testConfigure_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_279_elements(202) & testConfigure_CP_279_elements(203);
      gj_testConfigure_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_279_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  merge  transition  place  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	201 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_79/merge_stmt_363_PhiReqMerge
      -- CP-element group 205: 	 branch_block_stmt_79/merge_stmt_363_PhiAck/$entry
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(205)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(205)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(205) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_CP_279_elements(205) <= OrReduce(testConfigure_CP_279_elements(201) & testConfigure_CP_279_elements(204));
    -- CP-element group 206:  fork  transition  place  input  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	159 
    -- CP-element group 206: 	160 
    -- CP-element group 206:  members (11) 
      -- CP-element group 206: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_Update/ccr
      -- CP-element group 206: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_update_start_
      -- CP-element group 206: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/$entry
      -- CP-element group 206: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384/call_stmt_373_Sample/crr
      -- CP-element group 206: 	 branch_block_stmt_79/merge_stmt_363__exit__
      -- CP-element group 206: 	 branch_block_stmt_79/call_stmt_373_to_assign_stmt_384__entry__
      -- CP-element group 206: 	 branch_block_stmt_79/merge_stmt_363_PhiAck/$exit
      -- CP-element group 206: 	 branch_block_stmt_79/merge_stmt_363_PhiAck/phi_stmt_364_ack
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(206)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(206)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(206) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:phi_stmt_364_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:call_stmt_373_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:call_stmt_373_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_364_ack_1767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_364_ack_0, ack => testConfigure_CP_279_elements(206)); -- 
    ccr_1447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(206), ack => call_stmt_373_call_req_1); -- 
    crr_1442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_279_elements(206), ack => call_stmt_373_call_req_0); -- 
    -- CP-element group 207:  merge  transition  place  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	52 
    -- CP-element group 207: 	156 
    -- CP-element group 207: 	161 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (16) 
      -- CP-element group 207: 	 $exit
      -- CP-element group 207: 	 branch_block_stmt_79/$exit
      -- CP-element group 207: 	 branch_block_stmt_79/branch_block_stmt_79__exit__
      -- CP-element group 207: 	 branch_block_stmt_79/merge_stmt_393__exit__
      -- CP-element group 207: 	 branch_block_stmt_79/return__
      -- CP-element group 207: 	 branch_block_stmt_79/merge_stmt_395__exit__
      -- CP-element group 207: 	 branch_block_stmt_79/merge_stmt_393_PhiReqMerge
      -- CP-element group 207: 	 branch_block_stmt_79/merge_stmt_393_PhiAck/$entry
      -- CP-element group 207: 	 branch_block_stmt_79/merge_stmt_393_PhiAck/$exit
      -- CP-element group 207: 	 branch_block_stmt_79/merge_stmt_393_PhiAck/dummy
      -- CP-element group 207: 	 branch_block_stmt_79/return___PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_79/return___PhiReq/$exit
      -- CP-element group 207: 	 branch_block_stmt_79/merge_stmt_395_PhiReqMerge
      -- CP-element group 207: 	 branch_block_stmt_79/merge_stmt_395_PhiAck/$entry
      -- CP-element group 207: 	 branch_block_stmt_79/merge_stmt_395_PhiAck/$exit
      -- CP-element group 207: 	 branch_block_stmt_79/merge_stmt_395_PhiAck/dummy
      -- 
    -- logger for CP element group testConfigure_CP_279_elements(207)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and testConfigure_CP_279_elements(207)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:testConfigure:CP:testConfigure_CP_279_elements(207) fired."); 
        -- 
      end if; --
    end process; 
    testConfigure_CP_279_elements(207) <= OrReduce(testConfigure_CP_279_elements(52) & testConfigure_CP_279_elements(156) & testConfigure_CP_279_elements(161));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar65_165_resized : std_logic_vector(6 downto 0);
    signal R_indvar65_165_scaled : std_logic_vector(6 downto 0);
    signal R_indvar65_172_resized : std_logic_vector(8 downto 0);
    signal R_indvar65_172_scaled : std_logic_vector(8 downto 0);
    signal R_indvar_275_resized : std_logic_vector(8 downto 0);
    signal R_indvar_275_scaled : std_logic_vector(8 downto 0);
    signal array_obj_ref_166_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_166_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_166_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_166_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_166_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_166_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_173_constant_part_of_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_173_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_173_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_173_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_173_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_173_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_276_constant_part_of_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_276_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_276_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_276_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_276_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_276_root_address : std_logic_vector(8 downto 0);
    signal arrayidx21_278 : std_logic_vector(31 downto 0);
    signal arrayidx7_168 : std_logic_vector(31 downto 0);
    signal arrayidx_175 : std_logic_vector(31 downto 0);
    signal call3_189 : std_logic_vector(15 downto 0);
    signal call_178 : std_logic_vector(15 downto 0);
    signal cmp1648_136 : std_logic_vector(0 downto 0);
    signal cmp3445_324 : std_logic_vector(0 downto 0);
    signal cmp_218 : std_logic_vector(0 downto 0);
    signal conv4_193 : std_logic_vector(31 downto 0);
    signal conv_182 : std_logic_vector(31 downto 0);
    signal exitcond7_384 : std_logic_vector(0 downto 0);
    signal exitcond_298 : std_logic_vector(0 downto 0);
    signal iNsTr_0_85 : std_logic_vector(31 downto 0);
    signal iNsTr_13_209 : std_logic_vector(31 downto 0);
    signal iNsTr_17_241 : std_logic_vector(63 downto 0);
    signal iNsTr_22_364 : std_logic_vector(63 downto 0);
    signal iNsTr_2_96 : std_logic_vector(31 downto 0);
    signal iNsTr_4_107 : std_logic_vector(31 downto 0);
    signal iNsTr_6_118 : std_logic_vector(31 downto 0);
    signal inc_161 : std_logic_vector(31 downto 0);
    signal indvar65_144 : std_logic_vector(63 downto 0);
    signal indvar_257 : std_logic_vector(63 downto 0);
    signal indvarx_xnext58_293 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_379 : std_logic_vector(63 downto 0);
    signal mul_287 : std_logic_vector(31 downto 0);
    signal mulx_xlcssa_306 : std_logic_vector(31 downto 0);
    signal num_elemsx_x050_264 : std_logic_vector(31 downto 0);
    signal num_elemsx_x050x_xlcssa_314 : std_logic_vector(31 downto 0);
    signal ptr_deref_109_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_109_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_109_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_109_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_109_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_109_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_109_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_109_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_109_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_109_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_109_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_109_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_109_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_109_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_109_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_120_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_120_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_120_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_120_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_120_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_120_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_184_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_184_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_184_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_184_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_184_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_184_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_184_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_184_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_184_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_184_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_184_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_184_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_184_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_184_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_184_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_195_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_195_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_195_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_195_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_195_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_195_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_212_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_212_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_212_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_212_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_212_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_212_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_212_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_212_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_212_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_212_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_212_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_212_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_212_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_212_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_281_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_281_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_281_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_281_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_281_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_281_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_281_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_281_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_281_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_281_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_281_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_281_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_281_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_281_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_87_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_87_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_87_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_87_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_87_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_87_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_87_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_87_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_87_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_87_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_87_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_87_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_87_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_87_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_87_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_98_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_98_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_98_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_98_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_98_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_98_word_offset_0 : std_logic_vector(8 downto 0);
    signal tmp15x_xop_237 : std_logic_vector(31 downto 0);
    signal tmp1_213 : std_logic_vector(31 downto 0);
    signal tmp1x_xlcssa_126 : std_logic_vector(31 downto 0);
    signal tmp22_282 : std_logic_vector(31 downto 0);
    signal tmp22x_xlcssa_310 : std_logic_vector(31 downto 0);
    signal tmp2_336 : std_logic_vector(31 downto 0);
    signal tmp3_342 : std_logic_vector(63 downto 0);
    signal tmp4_348 : std_logic_vector(63 downto 0);
    signal tmp59_231 : std_logic_vector(0 downto 0);
    signal tmp5_354 : std_logic_vector(0 downto 0);
    signal tmp63_254 : std_logic_vector(63 downto 0);
    signal tmp67_203 : std_logic_vector(63 downto 0);
    signal tmp_157 : std_logic_vector(63 downto 0);
    signal type_cast_100_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_111_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_122_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_129_wire : std_logic_vector(31 downto 0);
    signal type_cast_134_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_148_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_150_wire : std_logic_vector(63 downto 0);
    signal type_cast_155_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_201_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_229_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_235_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_245_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_252_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_261_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_263_wire : std_logic_vector(63 downto 0);
    signal type_cast_268_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_270_wire : std_logic_vector(31 downto 0);
    signal type_cast_291_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_309_wire : std_logic_vector(31 downto 0);
    signal type_cast_313_wire : std_logic_vector(31 downto 0);
    signal type_cast_317_wire : std_logic_vector(31 downto 0);
    signal type_cast_322_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_340_wire : std_logic_vector(63 downto 0);
    signal type_cast_346_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_352_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_359_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_368_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_370_wire : std_logic_vector(63 downto 0);
    signal type_cast_377_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_89_wire_constant : std_logic_vector(31 downto 0);
    signal umax6_361 : std_logic_vector(63 downto 0);
    signal xx_xop_247 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_166_constant_part_of_offset <= "0000010";
    array_obj_ref_166_offset_scale_factor_0 <= "1000000";
    array_obj_ref_166_offset_scale_factor_1 <= "0000001";
    array_obj_ref_166_resized_base_address <= "0000000";
    array_obj_ref_173_constant_part_of_offset <= "000001001";
    array_obj_ref_173_offset_scale_factor_0 <= "100000000";
    array_obj_ref_173_offset_scale_factor_1 <= "000000100";
    array_obj_ref_173_resized_base_address <= "000000000";
    array_obj_ref_276_constant_part_of_offset <= "000001001";
    array_obj_ref_276_offset_scale_factor_0 <= "100000000";
    array_obj_ref_276_offset_scale_factor_1 <= "000000100";
    array_obj_ref_276_resized_base_address <= "000000000";
    iNsTr_0_85 <= "00000000000000000000000000000000";
    iNsTr_13_209 <= "00000000000000000000000000000101";
    iNsTr_2_96 <= "00000000000000000000000000000100";
    iNsTr_4_107 <= "00000000000000000000000000000101";
    iNsTr_6_118 <= "00000000000000000000000000000001";
    ptr_deref_109_word_offset_0 <= "000000000";
    ptr_deref_109_word_offset_1 <= "000000001";
    ptr_deref_109_word_offset_2 <= "000000010";
    ptr_deref_109_word_offset_3 <= "000000011";
    ptr_deref_120_word_offset_0 <= "0000000";
    ptr_deref_184_word_offset_0 <= "000000000";
    ptr_deref_184_word_offset_1 <= "000000001";
    ptr_deref_184_word_offset_2 <= "000000010";
    ptr_deref_184_word_offset_3 <= "000000011";
    ptr_deref_195_word_offset_0 <= "0000000";
    ptr_deref_212_word_offset_0 <= "000000000";
    ptr_deref_212_word_offset_1 <= "000000001";
    ptr_deref_212_word_offset_2 <= "000000010";
    ptr_deref_212_word_offset_3 <= "000000011";
    ptr_deref_281_word_offset_0 <= "000000000";
    ptr_deref_281_word_offset_1 <= "000000001";
    ptr_deref_281_word_offset_2 <= "000000010";
    ptr_deref_281_word_offset_3 <= "000000011";
    ptr_deref_87_word_offset_0 <= "000000000";
    ptr_deref_87_word_offset_1 <= "000000001";
    ptr_deref_87_word_offset_2 <= "000000010";
    ptr_deref_87_word_offset_3 <= "000000011";
    ptr_deref_98_word_offset_0 <= "000000000";
    type_cast_100_wire_constant <= "00000001";
    type_cast_111_wire_constant <= "00000000000000000000000000000011";
    type_cast_122_wire_constant <= "00000000000000000000000000000011";
    type_cast_134_wire_constant <= "00000000000000000000000000000000";
    type_cast_148_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_155_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_201_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_229_wire_constant <= "00000000000000000000000000000001";
    type_cast_235_wire_constant <= "11111111111111111111111111111111";
    type_cast_245_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_252_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_261_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_268_wire_constant <= "00000000000000000000000000000001";
    type_cast_291_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_322_wire_constant <= "00000000000000000000000000001111";
    type_cast_346_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_352_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_359_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_368_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_377_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_89_wire_constant <= "00000000000000000000000000000001";
    -- logger for phi phi_stmt_126
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_126_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_126:input-0 type_cast_129_wire= " & Convert_SLV_To_Hex_String(type_cast_129_wire));
          --
        end if;
        if phi_stmt_126_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:testConfigure:DP:phi_stmt_126:sample-completed");
          --
        end if;
        if phi_stmt_126_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:testConfigure:DP:phi_stmt_126:output tmp1x_xlcssa_126= " & Convert_SLV_To_Hex_String(tmp1x_xlcssa_126));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_126: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_129_wire;
      req(0) <= phi_stmt_126_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_126",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_126_ack_0,
          idata => idata,
          odata => tmp1x_xlcssa_126,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_126
    -- logger for phi phi_stmt_144
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_144_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_144:input-0 type_cast_148_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_148_wire_constant));
          --
        end if;
        if phi_stmt_144_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_144:input-1 type_cast_150_wire= " & Convert_SLV_To_Hex_String(type_cast_150_wire));
          --
        end if;
        if phi_stmt_144_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:testConfigure:DP:phi_stmt_144:sample-completed");
          --
        end if;
        if phi_stmt_144_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:testConfigure:DP:phi_stmt_144:output indvar65_144= " & Convert_SLV_To_Hex_String(indvar65_144));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_144: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_148_wire_constant & type_cast_150_wire;
      req <= phi_stmt_144_req_0 & phi_stmt_144_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_144",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_144_ack_0,
          idata => idata,
          odata => indvar65_144,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_144
    -- logger for phi phi_stmt_257
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_257_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_257:input-0 type_cast_261_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_261_wire_constant));
          --
        end if;
        if phi_stmt_257_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_257:input-1 type_cast_263_wire= " & Convert_SLV_To_Hex_String(type_cast_263_wire));
          --
        end if;
        if phi_stmt_257_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:testConfigure:DP:phi_stmt_257:sample-completed");
          --
        end if;
        if phi_stmt_257_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:testConfigure:DP:phi_stmt_257:output indvar_257= " & Convert_SLV_To_Hex_String(indvar_257));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_257: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_261_wire_constant & type_cast_263_wire;
      req <= phi_stmt_257_req_0 & phi_stmt_257_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_257",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_257_ack_0,
          idata => idata,
          odata => indvar_257,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_257
    -- logger for phi phi_stmt_264
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_264_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_264:input-0 type_cast_268_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_268_wire_constant));
          --
        end if;
        if phi_stmt_264_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_264:input-1 type_cast_270_wire= " & Convert_SLV_To_Hex_String(type_cast_270_wire));
          --
        end if;
        if phi_stmt_264_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:testConfigure:DP:phi_stmt_264:sample-completed");
          --
        end if;
        if phi_stmt_264_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:testConfigure:DP:phi_stmt_264:output num_elemsx_x050_264= " & Convert_SLV_To_Hex_String(num_elemsx_x050_264));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_264: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_268_wire_constant & type_cast_270_wire;
      req <= phi_stmt_264_req_0 & phi_stmt_264_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_264",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_264_ack_0,
          idata => idata,
          odata => num_elemsx_x050_264,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_264
    -- logger for phi phi_stmt_306
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_306_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_306:input-0 type_cast_309_wire= " & Convert_SLV_To_Hex_String(type_cast_309_wire));
          --
        end if;
        if phi_stmt_306_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:testConfigure:DP:phi_stmt_306:sample-completed");
          --
        end if;
        if phi_stmt_306_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:testConfigure:DP:phi_stmt_306:output mulx_xlcssa_306= " & Convert_SLV_To_Hex_String(mulx_xlcssa_306));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_306: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_309_wire;
      req(0) <= phi_stmt_306_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_306",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_306_ack_0,
          idata => idata,
          odata => mulx_xlcssa_306,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_306
    -- logger for phi phi_stmt_310
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_310_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_310:input-0 type_cast_313_wire= " & Convert_SLV_To_Hex_String(type_cast_313_wire));
          --
        end if;
        if phi_stmt_310_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:testConfigure:DP:phi_stmt_310:sample-completed");
          --
        end if;
        if phi_stmt_310_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:testConfigure:DP:phi_stmt_310:output tmp22x_xlcssa_310= " & Convert_SLV_To_Hex_String(tmp22x_xlcssa_310));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_310: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_313_wire;
      req(0) <= phi_stmt_310_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_310",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_310_ack_0,
          idata => idata,
          odata => tmp22x_xlcssa_310,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_310
    -- logger for phi phi_stmt_314
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_314_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_314:input-0 type_cast_317_wire= " & Convert_SLV_To_Hex_String(type_cast_317_wire));
          --
        end if;
        if phi_stmt_314_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:testConfigure:DP:phi_stmt_314:sample-completed");
          --
        end if;
        if phi_stmt_314_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:testConfigure:DP:phi_stmt_314:output num_elemsx_x050x_xlcssa_314= " & Convert_SLV_To_Hex_String(num_elemsx_x050x_xlcssa_314));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_314: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_317_wire;
      req(0) <= phi_stmt_314_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_314",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_314_ack_0,
          idata => idata,
          odata => num_elemsx_x050x_xlcssa_314,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_314
    -- logger for phi phi_stmt_364
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_364_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_364:input-0 type_cast_368_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_368_wire_constant));
          --
        end if;
        if phi_stmt_364_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:testConfigure:DP:phi_stmt_364:input-1 type_cast_370_wire= " & Convert_SLV_To_Hex_String(type_cast_370_wire));
          --
        end if;
        if phi_stmt_364_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:testConfigure:DP:phi_stmt_364:sample-completed");
          --
        end if;
        if phi_stmt_364_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:testConfigure:DP:phi_stmt_364:output iNsTr_22_364= " & Convert_SLV_To_Hex_String(iNsTr_22_364));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_364: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_368_wire_constant & type_cast_370_wire;
      req <= phi_stmt_364_req_0 & phi_stmt_364_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_364",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_364_ack_0,
          idata => idata,
          odata => iNsTr_22_364,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_364
    -- logger for split-operator MUX_253_inst flow-through 
    process(tmp63_254) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:MUX_253_inst:flowthrough inputs: " & " tmp59_231 = "& Convert_SLV_To_Hex_String(tmp59_231) & " xx_xop_247 = "& Convert_SLV_To_Hex_String(xx_xop_247) & " type_cast_252_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_252_wire_constant) & " outputs:" & " tmp63_254= "  & Convert_SLV_To_Hex_String(tmp63_254));
      --
    end process; 
    -- flow-through select operator MUX_253_inst
    tmp63_254 <= xx_xop_247 when (tmp59_231(0) /=  '0') else type_cast_252_wire_constant;
    -- logger for split-operator MUX_360_inst flow-through 
    process(umax6_361) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:MUX_360_inst:flowthrough inputs: " & " tmp5_354 = "& Convert_SLV_To_Hex_String(tmp5_354) & " tmp4_348 = "& Convert_SLV_To_Hex_String(tmp4_348) & " type_cast_359_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_359_wire_constant) & " outputs:" & " umax6_361= "  & Convert_SLV_To_Hex_String(umax6_361));
      --
    end process; 
    -- flow-through select operator MUX_360_inst
    umax6_361 <= tmp4_348 when (tmp5_354(0) /=  '0') else type_cast_359_wire_constant;
    -- logger for split-operator addr_of_167_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_167_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:addr_of_167_final_reg:started:   inputs: " & " array_obj_ref_166_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_166_root_address));
          --
        end if; 
        if addr_of_167_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:addr_of_167_final_reg:finished:  outputs: " & " arrayidx7_168= "  & Convert_SLV_To_Hex_String(arrayidx7_168));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_167_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_167_final_reg_req_0;
      addr_of_167_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_167_final_reg_req_1;
      addr_of_167_final_reg_ack_1<= rack(0);
      addr_of_167_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_167_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_166_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx7_168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_174_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_174_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:addr_of_174_final_reg:started:   inputs: " & " array_obj_ref_173_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_173_root_address));
          --
        end if; 
        if addr_of_174_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:addr_of_174_final_reg:finished:  outputs: " & " arrayidx_175= "  & Convert_SLV_To_Hex_String(arrayidx_175));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_174_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_174_final_reg_req_0;
      addr_of_174_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_174_final_reg_req_1;
      addr_of_174_final_reg_ack_1<= rack(0);
      addr_of_174_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_174_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 9,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_173_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator addr_of_277_final_reg
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if addr_of_277_final_reg_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:addr_of_277_final_reg:started:   inputs: " & " array_obj_ref_276_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_276_root_address));
          --
        end if; 
        if addr_of_277_final_reg_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:addr_of_277_final_reg:finished:  outputs: " & " arrayidx21_278= "  & Convert_SLV_To_Hex_String(arrayidx21_278));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    addr_of_277_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_277_final_reg_req_0;
      addr_of_277_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_277_final_reg_req_1;
      addr_of_277_final_reg_ack_1<= rack(0);
      addr_of_277_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_277_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 9,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_276_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx21_278,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_129_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_129_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_129_inst:started:   inputs: " & " tmp1_213 = "& Convert_SLV_To_Hex_String(tmp1_213));
          --
        end if; 
        if type_cast_129_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_129_inst:finished:  outputs: " & " type_cast_129_wire= "  & Convert_SLV_To_Hex_String(type_cast_129_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_129_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_129_inst_req_0;
      type_cast_129_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_129_inst_req_1;
      type_cast_129_inst_ack_1<= rack(0);
      type_cast_129_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_129_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_213,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_129_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_150_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_150_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_150_inst:started:   inputs: " & " tmp67_203 = "& Convert_SLV_To_Hex_String(tmp67_203));
          --
        end if; 
        if type_cast_150_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_150_inst:finished:  outputs: " & " type_cast_150_wire= "  & Convert_SLV_To_Hex_String(type_cast_150_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_150_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_150_inst_req_0;
      type_cast_150_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_150_inst_req_1;
      type_cast_150_inst_ack_1<= rack(0);
      type_cast_150_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_150_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp67_203,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_150_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_160_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_160_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_160_inst:started:   inputs: " & " tmp_157 = "& Convert_SLV_To_Hex_String(tmp_157));
          --
        end if; 
        if type_cast_160_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_160_inst:finished:  outputs: " & " inc_161= "  & Convert_SLV_To_Hex_String(inc_161));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_160_inst_req_0;
      type_cast_160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_160_inst_req_1;
      type_cast_160_inst_ack_1<= rack(0);
      type_cast_160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_181_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_181_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_181_inst:started:   inputs: " & " call_178 = "& Convert_SLV_To_Hex_String(call_178));
          --
        end if; 
        if type_cast_181_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_181_inst:finished:  outputs: " & " conv_182= "  & Convert_SLV_To_Hex_String(conv_182));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_181_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_181_inst_req_0;
      type_cast_181_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_181_inst_req_1;
      type_cast_181_inst_ack_1<= rack(0);
      type_cast_181_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_181_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_178,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_182,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_192_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_192_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_192_inst:started:   inputs: " & " call3_189 = "& Convert_SLV_To_Hex_String(call3_189));
          --
        end if; 
        if type_cast_192_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_192_inst:finished:  outputs: " & " conv4_193= "  & Convert_SLV_To_Hex_String(conv4_193));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_192_inst_req_0;
      type_cast_192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_192_inst_req_1;
      type_cast_192_inst_ack_1<= rack(0);
      type_cast_192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_189,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_240_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_240_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_240_inst:started:   inputs: " & " tmp15x_xop_237 = "& Convert_SLV_To_Hex_String(tmp15x_xop_237));
          --
        end if; 
        if type_cast_240_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_240_inst:finished:  outputs: " & " iNsTr_17_241= "  & Convert_SLV_To_Hex_String(iNsTr_17_241));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_240_inst_req_0;
      type_cast_240_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_240_inst_req_1;
      type_cast_240_inst_ack_1<= rack(0);
      type_cast_240_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_240_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp15x_xop_237,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_17_241,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_263_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_263_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_263_inst:started:   inputs: " & " indvarx_xnext58_293 = "& Convert_SLV_To_Hex_String(indvarx_xnext58_293));
          --
        end if; 
        if type_cast_263_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_263_inst:finished:  outputs: " & " type_cast_263_wire= "  & Convert_SLV_To_Hex_String(type_cast_263_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_263_inst_req_0;
      type_cast_263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_263_inst_req_1;
      type_cast_263_inst_ack_1<= rack(0);
      type_cast_263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext58_293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_263_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_270_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_270_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_270_inst:started:   inputs: " & " mul_287 = "& Convert_SLV_To_Hex_String(mul_287));
          --
        end if; 
        if type_cast_270_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_270_inst:finished:  outputs: " & " type_cast_270_wire= "  & Convert_SLV_To_Hex_String(type_cast_270_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_270_inst_req_0;
      type_cast_270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_270_inst_req_1;
      type_cast_270_inst_ack_1<= rack(0);
      type_cast_270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_270_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul_287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_270_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_309_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_309_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_309_inst:started:   inputs: " & " mul_287 = "& Convert_SLV_To_Hex_String(mul_287));
          --
        end if; 
        if type_cast_309_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_309_inst:finished:  outputs: " & " type_cast_309_wire= "  & Convert_SLV_To_Hex_String(type_cast_309_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_309_inst_req_0;
      type_cast_309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_309_inst_req_1;
      type_cast_309_inst_ack_1<= rack(0);
      type_cast_309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul_287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_309_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_313_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_313_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_313_inst:started:   inputs: " & " tmp22_282 = "& Convert_SLV_To_Hex_String(tmp22_282));
          --
        end if; 
        if type_cast_313_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_313_inst:finished:  outputs: " & " type_cast_313_wire= "  & Convert_SLV_To_Hex_String(type_cast_313_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_313_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_313_inst_req_0;
      type_cast_313_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_313_inst_req_1;
      type_cast_313_inst_ack_1<= rack(0);
      type_cast_313_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_313_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp22_282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_313_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_317_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_317_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_317_inst:started:   inputs: " & " num_elemsx_x050_264 = "& Convert_SLV_To_Hex_String(num_elemsx_x050_264));
          --
        end if; 
        if type_cast_317_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_317_inst:finished:  outputs: " & " type_cast_317_wire= "  & Convert_SLV_To_Hex_String(type_cast_317_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_317_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_317_inst_req_0;
      type_cast_317_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_317_inst_req_1;
      type_cast_317_inst_ack_1<= rack(0);
      type_cast_317_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_317_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_elemsx_x050_264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_317_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_341_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_341_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_341_inst:started:   inputs: " & " type_cast_340_wire = "& Convert_SLV_To_Hex_String(type_cast_340_wire));
          --
        end if; 
        if type_cast_341_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_341_inst:finished:  outputs: " & " tmp3_342= "  & Convert_SLV_To_Hex_String(tmp3_342));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_341_inst_req_0;
      type_cast_341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_341_inst_req_1;
      type_cast_341_inst_ack_1<= rack(0);
      type_cast_341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_340_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_370_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_370_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_370_inst:started:   inputs: " & " indvarx_xnext_379 = "& Convert_SLV_To_Hex_String(indvarx_xnext_379));
          --
        end if; 
        if type_cast_370_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_370_inst:finished:  outputs: " & " type_cast_370_wire= "  & Convert_SLV_To_Hex_String(type_cast_370_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_370_inst_req_0;
      type_cast_370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_370_inst_req_1;
      type_cast_370_inst_ack_1<= rack(0);
      type_cast_370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_379,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_370_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_166_index_1_rename flow-through 
    process(R_indvar65_165_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_166_index_1_rename:flowthrough  inputs: " & " R_indvar65_165_resized = "& Convert_SLV_To_Hex_String(R_indvar65_165_resized) & "outputs: " & " R_indvar65_165_scaled= "  & Convert_SLV_To_Hex_String(R_indvar65_165_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_166_index_1_rename
    process(R_indvar65_165_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar65_165_resized;
      ov(6 downto 0) := iv;
      R_indvar65_165_scaled <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_166_index_1_resize flow-through 
    process(R_indvar65_165_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_166_index_1_resize:flowthrough  inputs: " & " indvar65_144 = "& Convert_SLV_To_Hex_String(indvar65_144) & "outputs: " & " R_indvar65_165_resized= "  & Convert_SLV_To_Hex_String(R_indvar65_165_resized));
      --
    end process; 
    -- equivalence array_obj_ref_166_index_1_resize
    process(indvar65_144) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar65_144;
      ov := iv(6 downto 0);
      R_indvar65_165_resized <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_166_root_address_inst flow-through 
    process(array_obj_ref_166_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_166_root_address_inst:flowthrough  inputs: " & " array_obj_ref_166_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_166_final_offset) & "outputs: " & " array_obj_ref_166_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_166_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_166_root_address_inst
    process(array_obj_ref_166_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_166_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_166_root_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_173_index_1_resize flow-through 
    process(R_indvar65_172_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_173_index_1_resize:flowthrough  inputs: " & " indvar65_144 = "& Convert_SLV_To_Hex_String(indvar65_144) & "outputs: " & " R_indvar65_172_resized= "  & Convert_SLV_To_Hex_String(R_indvar65_172_resized));
      --
    end process; 
    -- equivalence array_obj_ref_173_index_1_resize
    process(indvar65_144) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar65_144;
      ov := iv(8 downto 0);
      R_indvar65_172_resized <= ov(8 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_173_root_address_inst flow-through 
    process(array_obj_ref_173_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_173_root_address_inst:flowthrough  inputs: " & " array_obj_ref_173_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_173_final_offset) & "outputs: " & " array_obj_ref_173_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_173_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_173_root_address_inst
    process(array_obj_ref_173_final_offset) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_173_final_offset;
      ov(8 downto 0) := iv;
      array_obj_ref_173_root_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_276_index_1_resize flow-through 
    process(R_indvar_275_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_276_index_1_resize:flowthrough  inputs: " & " indvar_257 = "& Convert_SLV_To_Hex_String(indvar_257) & "outputs: " & " R_indvar_275_resized= "  & Convert_SLV_To_Hex_String(R_indvar_275_resized));
      --
    end process; 
    -- equivalence array_obj_ref_276_index_1_resize
    process(indvar_257) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_257;
      ov := iv(8 downto 0);
      R_indvar_275_resized <= ov(8 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_276_root_address_inst flow-through 
    process(array_obj_ref_276_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_276_root_address_inst:flowthrough  inputs: " & " array_obj_ref_276_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_276_final_offset) & "outputs: " & " array_obj_ref_276_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_276_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_276_root_address_inst
    process(array_obj_ref_276_final_offset) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_276_final_offset;
      ov(8 downto 0) := iv;
      array_obj_ref_276_root_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_109_base_resize flow-through 
    process(ptr_deref_109_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_base_resize:flowthrough  inputs: " & " iNsTr_4_107 = "& Convert_SLV_To_Hex_String(iNsTr_4_107) & "outputs: " & " ptr_deref_109_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_109_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_109_base_resize
    process(iNsTr_4_107) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_107;
      ov := iv(8 downto 0);
      ptr_deref_109_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_109_gather_scatter flow-through 
    process(ptr_deref_109_data_3, ptr_deref_109_data_2, ptr_deref_109_data_1, ptr_deref_109_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_gather_scatter:flowthrough  inputs: " & " type_cast_111_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_111_wire_constant) & "outputs: " & " ptr_deref_109_data_3= "  & Convert_SLV_To_Hex_String(ptr_deref_109_data_3) & " ptr_deref_109_data_2= "  & Convert_SLV_To_Hex_String(ptr_deref_109_data_2) & " ptr_deref_109_data_1= "  & Convert_SLV_To_Hex_String(ptr_deref_109_data_1) & " ptr_deref_109_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_109_data_0));
      --
    end process; 
    -- equivalence ptr_deref_109_gather_scatter
    process(type_cast_111_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_111_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_109_data_3 <= ov(31 downto 24);
      ptr_deref_109_data_2 <= ov(23 downto 16);
      ptr_deref_109_data_1 <= ov(15 downto 8);
      ptr_deref_109_data_0 <= ov(7 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_109_root_address_inst flow-through 
    process(ptr_deref_109_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_root_address_inst:flowthrough  inputs: " & " ptr_deref_109_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_109_resized_base_address) & "outputs: " & " ptr_deref_109_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_109_root_address));
      --
    end process; 
    -- equivalence ptr_deref_109_root_address_inst
    process(ptr_deref_109_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_109_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_109_root_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_120_addr_0 flow-through 
    process(ptr_deref_120_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_120_addr_0:flowthrough  inputs: " & " ptr_deref_120_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_120_root_address) & "outputs: " & " ptr_deref_120_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_120_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_120_addr_0
    process(ptr_deref_120_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_120_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_120_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_120_base_resize flow-through 
    process(ptr_deref_120_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_120_base_resize:flowthrough  inputs: " & " iNsTr_6_118 = "& Convert_SLV_To_Hex_String(iNsTr_6_118) & "outputs: " & " ptr_deref_120_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_120_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_120_base_resize
    process(iNsTr_6_118) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_118;
      ov := iv(6 downto 0);
      ptr_deref_120_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_120_gather_scatter flow-through 
    process(ptr_deref_120_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_120_gather_scatter:flowthrough  inputs: " & " type_cast_122_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_122_wire_constant) & "outputs: " & " ptr_deref_120_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_120_data_0));
      --
    end process; 
    -- equivalence ptr_deref_120_gather_scatter
    process(type_cast_122_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_122_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_120_data_0 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_120_root_address_inst flow-through 
    process(ptr_deref_120_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_120_root_address_inst:flowthrough  inputs: " & " ptr_deref_120_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_120_resized_base_address) & "outputs: " & " ptr_deref_120_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_120_root_address));
      --
    end process; 
    -- equivalence ptr_deref_120_root_address_inst
    process(ptr_deref_120_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_120_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_120_root_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_184_base_resize flow-through 
    process(ptr_deref_184_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_base_resize:flowthrough  inputs: " & " arrayidx_175 = "& Convert_SLV_To_Hex_String(arrayidx_175) & "outputs: " & " ptr_deref_184_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_184_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_184_base_resize
    process(arrayidx_175) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_175;
      ov := iv(8 downto 0);
      ptr_deref_184_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_184_gather_scatter flow-through 
    process(ptr_deref_184_data_3, ptr_deref_184_data_2, ptr_deref_184_data_1, ptr_deref_184_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_gather_scatter:flowthrough  inputs: " & " conv_182 = "& Convert_SLV_To_Hex_String(conv_182) & "outputs: " & " ptr_deref_184_data_3= "  & Convert_SLV_To_Hex_String(ptr_deref_184_data_3) & " ptr_deref_184_data_2= "  & Convert_SLV_To_Hex_String(ptr_deref_184_data_2) & " ptr_deref_184_data_1= "  & Convert_SLV_To_Hex_String(ptr_deref_184_data_1) & " ptr_deref_184_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_184_data_0));
      --
    end process; 
    -- equivalence ptr_deref_184_gather_scatter
    process(conv_182) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_182;
      ov(31 downto 0) := iv;
      ptr_deref_184_data_3 <= ov(31 downto 24);
      ptr_deref_184_data_2 <= ov(23 downto 16);
      ptr_deref_184_data_1 <= ov(15 downto 8);
      ptr_deref_184_data_0 <= ov(7 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_184_root_address_inst flow-through 
    process(ptr_deref_184_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_root_address_inst:flowthrough  inputs: " & " ptr_deref_184_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_184_resized_base_address) & "outputs: " & " ptr_deref_184_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_184_root_address));
      --
    end process; 
    -- equivalence ptr_deref_184_root_address_inst
    process(ptr_deref_184_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_184_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_184_root_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_195_addr_0 flow-through 
    process(ptr_deref_195_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_195_addr_0:flowthrough  inputs: " & " ptr_deref_195_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_195_root_address) & "outputs: " & " ptr_deref_195_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_195_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_195_addr_0
    process(ptr_deref_195_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_195_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_195_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_195_base_resize flow-through 
    process(ptr_deref_195_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_195_base_resize:flowthrough  inputs: " & " arrayidx7_168 = "& Convert_SLV_To_Hex_String(arrayidx7_168) & "outputs: " & " ptr_deref_195_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_195_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_195_base_resize
    process(arrayidx7_168) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx7_168;
      ov := iv(6 downto 0);
      ptr_deref_195_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_195_gather_scatter flow-through 
    process(ptr_deref_195_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_195_gather_scatter:flowthrough  inputs: " & " conv4_193 = "& Convert_SLV_To_Hex_String(conv4_193) & "outputs: " & " ptr_deref_195_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_195_data_0));
      --
    end process; 
    -- equivalence ptr_deref_195_gather_scatter
    process(conv4_193) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4_193;
      ov(31 downto 0) := iv;
      ptr_deref_195_data_0 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_195_root_address_inst flow-through 
    process(ptr_deref_195_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_195_root_address_inst:flowthrough  inputs: " & " ptr_deref_195_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_195_resized_base_address) & "outputs: " & " ptr_deref_195_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_195_root_address));
      --
    end process; 
    -- equivalence ptr_deref_195_root_address_inst
    process(ptr_deref_195_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_195_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_195_root_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_212_base_resize flow-through 
    process(ptr_deref_212_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_base_resize:flowthrough  inputs: " & " iNsTr_13_209 = "& Convert_SLV_To_Hex_String(iNsTr_13_209) & "outputs: " & " ptr_deref_212_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_212_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_212_base_resize
    process(iNsTr_13_209) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_13_209;
      ov := iv(8 downto 0);
      ptr_deref_212_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_212_gather_scatter flow-through 
    process(tmp1_213) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_gather_scatter:flowthrough  inputs: " & " ptr_deref_212_data_3 = "& Convert_SLV_To_Hex_String(ptr_deref_212_data_3) & " ptr_deref_212_data_2 = "& Convert_SLV_To_Hex_String(ptr_deref_212_data_2) & " ptr_deref_212_data_1 = "& Convert_SLV_To_Hex_String(ptr_deref_212_data_1) & " ptr_deref_212_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_212_data_0) & "outputs: " & " tmp1_213= "  & Convert_SLV_To_Hex_String(tmp1_213));
      --
    end process; 
    -- equivalence ptr_deref_212_gather_scatter
    process(ptr_deref_212_data_3, ptr_deref_212_data_2, ptr_deref_212_data_1, ptr_deref_212_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_212_data_3 & ptr_deref_212_data_2 & ptr_deref_212_data_1 & ptr_deref_212_data_0;
      ov(31 downto 0) := iv;
      tmp1_213 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_212_root_address_inst flow-through 
    process(ptr_deref_212_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_root_address_inst:flowthrough  inputs: " & " ptr_deref_212_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_212_resized_base_address) & "outputs: " & " ptr_deref_212_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_212_root_address));
      --
    end process; 
    -- equivalence ptr_deref_212_root_address_inst
    process(ptr_deref_212_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_212_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_212_root_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_281_base_resize flow-through 
    process(ptr_deref_281_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_base_resize:flowthrough  inputs: " & " arrayidx21_278 = "& Convert_SLV_To_Hex_String(arrayidx21_278) & "outputs: " & " ptr_deref_281_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_281_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_281_base_resize
    process(arrayidx21_278) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx21_278;
      ov := iv(8 downto 0);
      ptr_deref_281_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_281_gather_scatter flow-through 
    process(tmp22_282) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_gather_scatter:flowthrough  inputs: " & " ptr_deref_281_data_3 = "& Convert_SLV_To_Hex_String(ptr_deref_281_data_3) & " ptr_deref_281_data_2 = "& Convert_SLV_To_Hex_String(ptr_deref_281_data_2) & " ptr_deref_281_data_1 = "& Convert_SLV_To_Hex_String(ptr_deref_281_data_1) & " ptr_deref_281_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_281_data_0) & "outputs: " & " tmp22_282= "  & Convert_SLV_To_Hex_String(tmp22_282));
      --
    end process; 
    -- equivalence ptr_deref_281_gather_scatter
    process(ptr_deref_281_data_3, ptr_deref_281_data_2, ptr_deref_281_data_1, ptr_deref_281_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_281_data_3 & ptr_deref_281_data_2 & ptr_deref_281_data_1 & ptr_deref_281_data_0;
      ov(31 downto 0) := iv;
      tmp22_282 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_281_root_address_inst flow-through 
    process(ptr_deref_281_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_root_address_inst:flowthrough  inputs: " & " ptr_deref_281_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_281_resized_base_address) & "outputs: " & " ptr_deref_281_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_281_root_address));
      --
    end process; 
    -- equivalence ptr_deref_281_root_address_inst
    process(ptr_deref_281_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_281_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_281_root_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_87_base_resize flow-through 
    process(ptr_deref_87_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_base_resize:flowthrough  inputs: " & " iNsTr_0_85 = "& Convert_SLV_To_Hex_String(iNsTr_0_85) & "outputs: " & " ptr_deref_87_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_87_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_87_base_resize
    process(iNsTr_0_85) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_85;
      ov := iv(8 downto 0);
      ptr_deref_87_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_87_gather_scatter flow-through 
    process(ptr_deref_87_data_3, ptr_deref_87_data_2, ptr_deref_87_data_1, ptr_deref_87_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_gather_scatter:flowthrough  inputs: " & " type_cast_89_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_89_wire_constant) & "outputs: " & " ptr_deref_87_data_3= "  & Convert_SLV_To_Hex_String(ptr_deref_87_data_3) & " ptr_deref_87_data_2= "  & Convert_SLV_To_Hex_String(ptr_deref_87_data_2) & " ptr_deref_87_data_1= "  & Convert_SLV_To_Hex_String(ptr_deref_87_data_1) & " ptr_deref_87_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_87_data_0));
      --
    end process; 
    -- equivalence ptr_deref_87_gather_scatter
    process(type_cast_89_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_89_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_87_data_3 <= ov(31 downto 24);
      ptr_deref_87_data_2 <= ov(23 downto 16);
      ptr_deref_87_data_1 <= ov(15 downto 8);
      ptr_deref_87_data_0 <= ov(7 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_87_root_address_inst flow-through 
    process(ptr_deref_87_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_root_address_inst:flowthrough  inputs: " & " ptr_deref_87_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_87_resized_base_address) & "outputs: " & " ptr_deref_87_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_87_root_address));
      --
    end process; 
    -- equivalence ptr_deref_87_root_address_inst
    process(ptr_deref_87_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_87_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_87_root_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_98_addr_0 flow-through 
    process(ptr_deref_98_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_98_addr_0:flowthrough  inputs: " & " ptr_deref_98_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_98_root_address) & "outputs: " & " ptr_deref_98_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_98_word_address_0));
      --
    end process; 
    -- equivalence ptr_deref_98_addr_0
    process(ptr_deref_98_root_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_98_root_address;
      ov(8 downto 0) := iv;
      ptr_deref_98_word_address_0 <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_98_base_resize flow-through 
    process(ptr_deref_98_resized_base_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_98_base_resize:flowthrough  inputs: " & " iNsTr_2_96 = "& Convert_SLV_To_Hex_String(iNsTr_2_96) & "outputs: " & " ptr_deref_98_resized_base_address= "  & Convert_SLV_To_Hex_String(ptr_deref_98_resized_base_address));
      --
    end process; 
    -- equivalence ptr_deref_98_base_resize
    process(iNsTr_2_96) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_96;
      ov := iv(8 downto 0);
      ptr_deref_98_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_98_gather_scatter flow-through 
    process(ptr_deref_98_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_98_gather_scatter:flowthrough  inputs: " & " type_cast_100_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_100_wire_constant) & "outputs: " & " ptr_deref_98_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_98_data_0));
      --
    end process; 
    -- equivalence ptr_deref_98_gather_scatter
    process(type_cast_100_wire_constant) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_100_wire_constant;
      ov(7 downto 0) := iv;
      ptr_deref_98_data_0 <= ov(7 downto 0);
      --
    end process;
    -- logger for operator ptr_deref_98_root_address_inst flow-through 
    process(ptr_deref_98_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_98_root_address_inst:flowthrough  inputs: " & " ptr_deref_98_resized_base_address = "& Convert_SLV_To_Hex_String(ptr_deref_98_resized_base_address) & "outputs: " & " ptr_deref_98_root_address= "  & Convert_SLV_To_Hex_String(ptr_deref_98_root_address));
      --
    end process; 
    -- equivalence ptr_deref_98_root_address_inst
    process(ptr_deref_98_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_98_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_98_root_address <= ov(8 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_137_branch_req_0," req0 if_stmt_137_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_137_branch_ack_0," ack0 if_stmt_137_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_137_branch_ack_1," ack1 if_stmt_137_branch");
    if_stmt_137_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1648_136;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_137_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_137_branch_req_0,
          ack0 => if_stmt_137_branch_ack_0,
          ack1 => if_stmt_137_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_219_branch_req_0," req0 if_stmt_219_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_219_branch_ack_0," ack0 if_stmt_219_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_219_branch_ack_1," ack1 if_stmt_219_branch");
    if_stmt_219_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_218;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_219_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_219_branch_req_0,
          ack0 => if_stmt_219_branch_ack_0,
          ack1 => if_stmt_219_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_299_branch_req_0," req0 if_stmt_299_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_299_branch_ack_0," ack0 if_stmt_299_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_299_branch_ack_1," ack1 if_stmt_299_branch");
    if_stmt_299_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_298;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_299_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_299_branch_req_0,
          ack0 => if_stmt_299_branch_ack_0,
          ack1 => if_stmt_299_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_325_branch_req_0," req0 if_stmt_325_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_325_branch_ack_0," ack0 if_stmt_325_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_325_branch_ack_1," ack1 if_stmt_325_branch");
    if_stmt_325_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp3445_324;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_325_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_325_branch_req_0,
          ack0 => if_stmt_325_branch_ack_0,
          ack1 => if_stmt_325_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_385_branch_req_0," req0 if_stmt_385_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_385_branch_ack_0," ack0 if_stmt_385_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_385_branch_ack_1," ack1 if_stmt_385_branch");
    if_stmt_385_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond7_384;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_385_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_385_branch_req_0,
          ack0 => if_stmt_385_branch_ack_0,
          ack1 => if_stmt_385_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u32_u32_236_inst flow-through 
    process(tmp15x_xop_237) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ADD_u32_u32_236_inst:flowthrough inputs: " & " tmp1x_xlcssa_126 = "& Convert_SLV_To_Hex_String(tmp1x_xlcssa_126) & " type_cast_235_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_235_wire_constant) & " outputs:" & " tmp15x_xop_237= "  & Convert_SLV_To_Hex_String(tmp15x_xop_237));
      --
    end process; 
    -- binary operator ADD_u32_u32_236_inst
    process(tmp1x_xlcssa_126) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1x_xlcssa_126, type_cast_235_wire_constant, tmp_var);
      tmp15x_xop_237 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_156_inst flow-through 
    process(tmp_157) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ADD_u64_u64_156_inst:flowthrough inputs: " & " indvar65_144 = "& Convert_SLV_To_Hex_String(indvar65_144) & " type_cast_155_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_155_wire_constant) & " outputs:" & " tmp_157= "  & Convert_SLV_To_Hex_String(tmp_157));
      --
    end process; 
    -- binary operator ADD_u64_u64_156_inst
    process(indvar65_144) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar65_144, type_cast_155_wire_constant, tmp_var);
      tmp_157 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_202_inst flow-through 
    process(tmp67_203) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ADD_u64_u64_202_inst:flowthrough inputs: " & " indvar65_144 = "& Convert_SLV_To_Hex_String(indvar65_144) & " type_cast_201_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_201_wire_constant) & " outputs:" & " tmp67_203= "  & Convert_SLV_To_Hex_String(tmp67_203));
      --
    end process; 
    -- binary operator ADD_u64_u64_202_inst
    process(indvar65_144) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar65_144, type_cast_201_wire_constant, tmp_var);
      tmp67_203 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_246_inst flow-through 
    process(xx_xop_247) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ADD_u64_u64_246_inst:flowthrough inputs: " & " iNsTr_17_241 = "& Convert_SLV_To_Hex_String(iNsTr_17_241) & " type_cast_245_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_245_wire_constant) & " outputs:" & " xx_xop_247= "  & Convert_SLV_To_Hex_String(xx_xop_247));
      --
    end process; 
    -- binary operator ADD_u64_u64_246_inst
    process(iNsTr_17_241) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_17_241, type_cast_245_wire_constant, tmp_var);
      xx_xop_247 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_292_inst flow-through 
    process(indvarx_xnext58_293) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ADD_u64_u64_292_inst:flowthrough inputs: " & " indvar_257 = "& Convert_SLV_To_Hex_String(indvar_257) & " type_cast_291_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_291_wire_constant) & " outputs:" & " indvarx_xnext58_293= "  & Convert_SLV_To_Hex_String(indvarx_xnext58_293));
      --
    end process; 
    -- binary operator ADD_u64_u64_292_inst
    process(indvar_257) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_257, type_cast_291_wire_constant, tmp_var);
      indvarx_xnext58_293 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u64_u64_378_inst flow-through 
    process(indvarx_xnext_379) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ADD_u64_u64_378_inst:flowthrough inputs: " & " iNsTr_22_364 = "& Convert_SLV_To_Hex_String(iNsTr_22_364) & " type_cast_377_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_377_wire_constant) & " outputs:" & " indvarx_xnext_379= "  & Convert_SLV_To_Hex_String(indvarx_xnext_379));
      --
    end process; 
    -- binary operator ADD_u64_u64_378_inst
    process(iNsTr_22_364) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_22_364, type_cast_377_wire_constant, tmp_var);
      indvarx_xnext_379 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u32_u1_135_inst flow-through 
    process(cmp1648_136) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:EQ_u32_u1_135_inst:flowthrough inputs: " & " tmp1x_xlcssa_126 = "& Convert_SLV_To_Hex_String(tmp1x_xlcssa_126) & " type_cast_134_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_134_wire_constant) & " outputs:" & " cmp1648_136= "  & Convert_SLV_To_Hex_String(cmp1648_136));
      --
    end process; 
    -- binary operator EQ_u32_u1_135_inst
    process(tmp1x_xlcssa_126) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tmp1x_xlcssa_126, type_cast_134_wire_constant, tmp_var);
      cmp1648_136 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_297_inst flow-through 
    process(exitcond_298) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:EQ_u64_u1_297_inst:flowthrough inputs: " & " indvarx_xnext58_293 = "& Convert_SLV_To_Hex_String(indvarx_xnext58_293) & " tmp63_254 = "& Convert_SLV_To_Hex_String(tmp63_254) & " outputs:" & " exitcond_298= "  & Convert_SLV_To_Hex_String(exitcond_298));
      --
    end process; 
    -- binary operator EQ_u64_u1_297_inst
    process(indvarx_xnext58_293, tmp63_254) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext58_293, tmp63_254, tmp_var);
      exitcond_298 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_383_inst flow-through 
    process(exitcond7_384) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:EQ_u64_u1_383_inst:flowthrough inputs: " & " indvarx_xnext_379 = "& Convert_SLV_To_Hex_String(indvarx_xnext_379) & " umax6_361 = "& Convert_SLV_To_Hex_String(umax6_361) & " outputs:" & " exitcond7_384= "  & Convert_SLV_To_Hex_String(exitcond7_384));
      --
    end process; 
    -- binary operator EQ_u64_u1_383_inst
    process(indvarx_xnext_379, umax6_361) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_379, umax6_361, tmp_var);
      exitcond7_384 <= tmp_var; --
    end process;
    -- logger for split-operator LSHR_u64_u64_347_inst flow-through 
    process(tmp4_348) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:LSHR_u64_u64_347_inst:flowthrough inputs: " & " tmp3_342 = "& Convert_SLV_To_Hex_String(tmp3_342) & " type_cast_346_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_346_wire_constant) & " outputs:" & " tmp4_348= "  & Convert_SLV_To_Hex_String(tmp4_348));
      --
    end process; 
    -- binary operator LSHR_u64_u64_347_inst
    process(tmp3_342) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp3_342, type_cast_346_wire_constant, tmp_var);
      tmp4_348 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_286_inst flow-through 
    process(mul_287) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:MUL_u32_u32_286_inst:flowthrough inputs: " & " tmp22_282 = "& Convert_SLV_To_Hex_String(tmp22_282) & " num_elemsx_x050_264 = "& Convert_SLV_To_Hex_String(num_elemsx_x050_264) & " outputs:" & " mul_287= "  & Convert_SLV_To_Hex_String(mul_287));
      --
    end process; 
    -- binary operator MUL_u32_u32_286_inst
    process(tmp22_282, num_elemsx_x050_264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp22_282, num_elemsx_x050_264, tmp_var);
      mul_287 <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u32_u32_335_inst flow-through 
    process(tmp2_336) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:MUL_u32_u32_335_inst:flowthrough inputs: " & " num_elemsx_x050x_xlcssa_314 = "& Convert_SLV_To_Hex_String(num_elemsx_x050x_xlcssa_314) & " tmp22x_xlcssa_310 = "& Convert_SLV_To_Hex_String(tmp22x_xlcssa_310) & " outputs:" & " tmp2_336= "  & Convert_SLV_To_Hex_String(tmp2_336));
      --
    end process; 
    -- binary operator MUL_u32_u32_335_inst
    process(num_elemsx_x050x_xlcssa_314, tmp22x_xlcssa_310) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(num_elemsx_x050x_xlcssa_314, tmp22x_xlcssa_310, tmp_var);
      tmp2_336 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u32_u1_230_inst flow-through 
    process(tmp59_231) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:UGT_u32_u1_230_inst:flowthrough inputs: " & " tmp1x_xlcssa_126 = "& Convert_SLV_To_Hex_String(tmp1x_xlcssa_126) & " type_cast_229_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_229_wire_constant) & " outputs:" & " tmp59_231= "  & Convert_SLV_To_Hex_String(tmp59_231));
      --
    end process; 
    -- binary operator UGT_u32_u1_230_inst
    process(tmp1x_xlcssa_126) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp1x_xlcssa_126, type_cast_229_wire_constant, tmp_var);
      tmp59_231 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u32_u1_323_inst flow-through 
    process(cmp3445_324) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:UGT_u32_u1_323_inst:flowthrough inputs: " & " mulx_xlcssa_306 = "& Convert_SLV_To_Hex_String(mulx_xlcssa_306) & " type_cast_322_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_322_wire_constant) & " outputs:" & " cmp3445_324= "  & Convert_SLV_To_Hex_String(cmp3445_324));
      --
    end process; 
    -- binary operator UGT_u32_u1_323_inst
    process(mulx_xlcssa_306) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mulx_xlcssa_306, type_cast_322_wire_constant, tmp_var);
      cmp3445_324 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u64_u1_353_inst flow-through 
    process(tmp5_354) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:UGT_u64_u1_353_inst:flowthrough inputs: " & " tmp4_348 = "& Convert_SLV_To_Hex_String(tmp4_348) & " type_cast_352_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_352_wire_constant) & " outputs:" & " tmp5_354= "  & Convert_SLV_To_Hex_String(tmp5_354));
      --
    end process; 
    -- binary operator UGT_u64_u1_353_inst
    process(tmp4_348) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp4_348, type_cast_352_wire_constant, tmp_var);
      tmp5_354 <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u32_u1_217_inst flow-through 
    process(cmp_218) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ULT_u32_u1_217_inst:flowthrough inputs: " & " inc_161 = "& Convert_SLV_To_Hex_String(inc_161) & " tmp1_213 = "& Convert_SLV_To_Hex_String(tmp1_213) & " outputs:" & " cmp_218= "  & Convert_SLV_To_Hex_String(cmp_218));
      --
    end process; 
    -- binary operator ULT_u32_u1_217_inst
    process(inc_161, tmp1_213) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc_161, tmp1_213, tmp_var);
      cmp_218 <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_166_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_166_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_166_index_offset:started:   inputs: " & " R_indvar65_165_scaled = "& Convert_SLV_To_Hex_String(R_indvar65_165_scaled) & " array_obj_ref_166_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_166_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_166_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_166_index_offset:finished:  outputs: " & " array_obj_ref_166_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_166_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (16) : array_obj_ref_166_index_offset 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar65_165_scaled;
      array_obj_ref_166_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_166_index_offset_req_0;
      array_obj_ref_166_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_166_index_offset_req_1;
      array_obj_ref_166_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000010",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- logger for split-operator array_obj_ref_276_index_1_scale
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_276_index_1_scale_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_276_index_1_scale:started:   inputs: " & " R_indvar_275_resized = "& Convert_SLV_To_Hex_String(R_indvar_275_resized) & " array_obj_ref_276_offset_scale_factor_1 = "& Convert_SLV_To_Hex_String(array_obj_ref_276_offset_scale_factor_1));
          --
        end if; 
        if array_obj_ref_276_index_1_scale_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_276_index_1_scale:finished:  outputs: " & " R_indvar_275_scaled= "  & Convert_SLV_To_Hex_String(R_indvar_275_scaled));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_173_index_1_scale
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_173_index_1_scale_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_173_index_1_scale:started:   inputs: " & " R_indvar65_172_resized = "& Convert_SLV_To_Hex_String(R_indvar65_172_resized) & " array_obj_ref_173_offset_scale_factor_1 = "& Convert_SLV_To_Hex_String(array_obj_ref_173_offset_scale_factor_1));
          --
        end if; 
        if array_obj_ref_173_index_1_scale_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_173_index_1_scale:finished:  outputs: " & " R_indvar65_172_scaled= "  & Convert_SLV_To_Hex_String(R_indvar65_172_scaled));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (17) : array_obj_ref_276_index_1_scale array_obj_ref_173_index_1_scale 
    ApIntMul_group_17: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(17 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_275_resized & R_indvar65_172_resized;
      R_indvar_275_scaled <= data_out(17 downto 9);
      R_indvar65_172_scaled <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      reqL_unguarded(1) <= array_obj_ref_276_index_1_scale_req_0;
      reqL_unguarded(0) <= array_obj_ref_173_index_1_scale_req_0;
      array_obj_ref_276_index_1_scale_ack_0 <= ackL_unguarded(1);
      array_obj_ref_173_index_1_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= array_obj_ref_276_index_1_scale_req_1;
      reqR_unguarded(0) <= array_obj_ref_173_index_1_scale_req_1;
      array_obj_ref_276_index_1_scale_ack_1 <= ackR_unguarded(1);
      array_obj_ref_173_index_1_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_17_accessRegulator_0: access_regulator_base generic map (name => "ApIntMul_group_17_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApIntMul_group_17_accessRegulator_1: access_regulator_base generic map (name => "ApIntMul_group_17_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApIntMul_group_17_gI: SplitGuardInterface generic map(name => "ApIntMul_group_17_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          name => "ApIntMul_group_17",
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000100",
          constant_width => 9,
          use_constant  => true,
          full_rate  => false,
          no_arbitration => false,
          min_clock_period => false,
          num_reqs => 2,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs --
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- logger for split-operator array_obj_ref_173_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_173_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_173_index_offset:started:   inputs: " & " R_indvar65_172_scaled = "& Convert_SLV_To_Hex_String(R_indvar65_172_scaled) & " array_obj_ref_173_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_173_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_173_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_173_index_offset:finished:  outputs: " & " array_obj_ref_173_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_173_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (18) : array_obj_ref_173_index_offset 
    ApIntAdd_group_18: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar65_172_scaled;
      array_obj_ref_173_final_offset <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_173_index_offset_req_0;
      array_obj_ref_173_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_173_index_offset_req_1;
      array_obj_ref_173_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_18_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_18_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_18",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000001001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- logger for split-operator array_obj_ref_276_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_276_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_276_index_offset:started:   inputs: " & " R_indvar_275_scaled = "& Convert_SLV_To_Hex_String(R_indvar_275_scaled) & " array_obj_ref_276_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_276_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_276_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:array_obj_ref_276_index_offset:finished:  outputs: " & " array_obj_ref_276_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_276_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (19) : array_obj_ref_276_index_offset 
    ApIntAdd_group_19: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_275_scaled;
      array_obj_ref_276_final_offset <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_276_index_offset_req_0;
      array_obj_ref_276_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_276_index_offset_req_1;
      array_obj_ref_276_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_19_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_19_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_19",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000001001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- logger for split-operator ptr_deref_109_addr_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_109_addr_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_addr_0:started:   inputs: " & " ptr_deref_109_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_109_root_address) & " ptr_deref_109_word_offset_0 = "& Convert_SLV_To_Hex_String(ptr_deref_109_word_offset_0));
          --
        end if; 
        if ptr_deref_109_addr_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_addr_0:finished:  outputs: " & " ptr_deref_109_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_109_word_address_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (20) : ptr_deref_109_addr_0 
    ApIntAdd_group_20: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_109_root_address;
      ptr_deref_109_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_109_addr_0_req_0;
      ptr_deref_109_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_109_addr_0_req_1;
      ptr_deref_109_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_20_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_20_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_20",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- logger for split-operator ptr_deref_109_addr_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_109_addr_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_addr_1:started:   inputs: " & " ptr_deref_109_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_109_root_address) & " ptr_deref_109_word_offset_1 = "& Convert_SLV_To_Hex_String(ptr_deref_109_word_offset_1));
          --
        end if; 
        if ptr_deref_109_addr_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_addr_1:finished:  outputs: " & " ptr_deref_109_word_address_1= "  & Convert_SLV_To_Hex_String(ptr_deref_109_word_address_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (21) : ptr_deref_109_addr_1 
    ApIntAdd_group_21: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_109_root_address;
      ptr_deref_109_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_109_addr_1_req_0;
      ptr_deref_109_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_109_addr_1_req_1;
      ptr_deref_109_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_21_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_21_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_21",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- logger for split-operator ptr_deref_109_addr_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_109_addr_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_addr_2:started:   inputs: " & " ptr_deref_109_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_109_root_address) & " ptr_deref_109_word_offset_2 = "& Convert_SLV_To_Hex_String(ptr_deref_109_word_offset_2));
          --
        end if; 
        if ptr_deref_109_addr_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_addr_2:finished:  outputs: " & " ptr_deref_109_word_address_2= "  & Convert_SLV_To_Hex_String(ptr_deref_109_word_address_2));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (22) : ptr_deref_109_addr_2 
    ApIntAdd_group_22: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_109_root_address;
      ptr_deref_109_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_109_addr_2_req_0;
      ptr_deref_109_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_109_addr_2_req_1;
      ptr_deref_109_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_22_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_22_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_22",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- logger for split-operator ptr_deref_109_addr_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_109_addr_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_addr_3:started:   inputs: " & " ptr_deref_109_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_109_root_address) & " ptr_deref_109_word_offset_3 = "& Convert_SLV_To_Hex_String(ptr_deref_109_word_offset_3));
          --
        end if; 
        if ptr_deref_109_addr_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_addr_3:finished:  outputs: " & " ptr_deref_109_word_address_3= "  & Convert_SLV_To_Hex_String(ptr_deref_109_word_address_3));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (23) : ptr_deref_109_addr_3 
    ApIntAdd_group_23: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_109_root_address;
      ptr_deref_109_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_109_addr_3_req_0;
      ptr_deref_109_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_109_addr_3_req_1;
      ptr_deref_109_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_23_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- logger for split-operator ptr_deref_184_addr_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_184_addr_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_addr_0:started:   inputs: " & " ptr_deref_184_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_184_root_address) & " ptr_deref_184_word_offset_0 = "& Convert_SLV_To_Hex_String(ptr_deref_184_word_offset_0));
          --
        end if; 
        if ptr_deref_184_addr_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_addr_0:finished:  outputs: " & " ptr_deref_184_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_184_word_address_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (24) : ptr_deref_184_addr_0 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_184_root_address;
      ptr_deref_184_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_184_addr_0_req_0;
      ptr_deref_184_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_184_addr_0_req_1;
      ptr_deref_184_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_24_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- logger for split-operator ptr_deref_184_addr_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_184_addr_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_addr_1:started:   inputs: " & " ptr_deref_184_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_184_root_address) & " ptr_deref_184_word_offset_1 = "& Convert_SLV_To_Hex_String(ptr_deref_184_word_offset_1));
          --
        end if; 
        if ptr_deref_184_addr_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_addr_1:finished:  outputs: " & " ptr_deref_184_word_address_1= "  & Convert_SLV_To_Hex_String(ptr_deref_184_word_address_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (25) : ptr_deref_184_addr_1 
    ApIntAdd_group_25: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_184_root_address;
      ptr_deref_184_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_184_addr_1_req_0;
      ptr_deref_184_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_184_addr_1_req_1;
      ptr_deref_184_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_25_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_25_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_25",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- logger for split-operator ptr_deref_184_addr_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_184_addr_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_addr_2:started:   inputs: " & " ptr_deref_184_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_184_root_address) & " ptr_deref_184_word_offset_2 = "& Convert_SLV_To_Hex_String(ptr_deref_184_word_offset_2));
          --
        end if; 
        if ptr_deref_184_addr_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_addr_2:finished:  outputs: " & " ptr_deref_184_word_address_2= "  & Convert_SLV_To_Hex_String(ptr_deref_184_word_address_2));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (26) : ptr_deref_184_addr_2 
    ApIntAdd_group_26: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_184_root_address;
      ptr_deref_184_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_184_addr_2_req_0;
      ptr_deref_184_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_184_addr_2_req_1;
      ptr_deref_184_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_26_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_26_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_26",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- logger for split-operator ptr_deref_184_addr_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_184_addr_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_addr_3:started:   inputs: " & " ptr_deref_184_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_184_root_address) & " ptr_deref_184_word_offset_3 = "& Convert_SLV_To_Hex_String(ptr_deref_184_word_offset_3));
          --
        end if; 
        if ptr_deref_184_addr_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_addr_3:finished:  outputs: " & " ptr_deref_184_word_address_3= "  & Convert_SLV_To_Hex_String(ptr_deref_184_word_address_3));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (27) : ptr_deref_184_addr_3 
    ApIntAdd_group_27: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_184_root_address;
      ptr_deref_184_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_184_addr_3_req_0;
      ptr_deref_184_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_184_addr_3_req_1;
      ptr_deref_184_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_27_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_27_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- logger for split-operator ptr_deref_212_addr_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_212_addr_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_addr_0:started:   inputs: " & " ptr_deref_212_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_212_root_address) & " ptr_deref_212_word_offset_0 = "& Convert_SLV_To_Hex_String(ptr_deref_212_word_offset_0));
          --
        end if; 
        if ptr_deref_212_addr_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_addr_0:finished:  outputs: " & " ptr_deref_212_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_212_word_address_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (28) : ptr_deref_212_addr_0 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_212_root_address;
      ptr_deref_212_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_212_addr_0_req_0;
      ptr_deref_212_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_212_addr_0_req_1;
      ptr_deref_212_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- logger for split-operator ptr_deref_212_addr_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_212_addr_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_addr_1:started:   inputs: " & " ptr_deref_212_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_212_root_address) & " ptr_deref_212_word_offset_1 = "& Convert_SLV_To_Hex_String(ptr_deref_212_word_offset_1));
          --
        end if; 
        if ptr_deref_212_addr_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_addr_1:finished:  outputs: " & " ptr_deref_212_word_address_1= "  & Convert_SLV_To_Hex_String(ptr_deref_212_word_address_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (29) : ptr_deref_212_addr_1 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_212_root_address;
      ptr_deref_212_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_212_addr_1_req_0;
      ptr_deref_212_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_212_addr_1_req_1;
      ptr_deref_212_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- logger for split-operator ptr_deref_212_addr_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_212_addr_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_addr_2:started:   inputs: " & " ptr_deref_212_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_212_root_address) & " ptr_deref_212_word_offset_2 = "& Convert_SLV_To_Hex_String(ptr_deref_212_word_offset_2));
          --
        end if; 
        if ptr_deref_212_addr_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_addr_2:finished:  outputs: " & " ptr_deref_212_word_address_2= "  & Convert_SLV_To_Hex_String(ptr_deref_212_word_address_2));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (30) : ptr_deref_212_addr_2 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_212_root_address;
      ptr_deref_212_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_212_addr_2_req_0;
      ptr_deref_212_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_212_addr_2_req_1;
      ptr_deref_212_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- logger for split-operator ptr_deref_212_addr_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_212_addr_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_addr_3:started:   inputs: " & " ptr_deref_212_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_212_root_address) & " ptr_deref_212_word_offset_3 = "& Convert_SLV_To_Hex_String(ptr_deref_212_word_offset_3));
          --
        end if; 
        if ptr_deref_212_addr_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_addr_3:finished:  outputs: " & " ptr_deref_212_word_address_3= "  & Convert_SLV_To_Hex_String(ptr_deref_212_word_address_3));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (31) : ptr_deref_212_addr_3 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_212_root_address;
      ptr_deref_212_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_212_addr_3_req_0;
      ptr_deref_212_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_212_addr_3_req_1;
      ptr_deref_212_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- logger for split-operator ptr_deref_281_addr_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_281_addr_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_addr_0:started:   inputs: " & " ptr_deref_281_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_281_root_address) & " ptr_deref_281_word_offset_0 = "& Convert_SLV_To_Hex_String(ptr_deref_281_word_offset_0));
          --
        end if; 
        if ptr_deref_281_addr_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_addr_0:finished:  outputs: " & " ptr_deref_281_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_281_word_address_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (32) : ptr_deref_281_addr_0 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_281_root_address;
      ptr_deref_281_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_281_addr_0_req_0;
      ptr_deref_281_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_281_addr_0_req_1;
      ptr_deref_281_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- logger for split-operator ptr_deref_281_addr_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_281_addr_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_addr_1:started:   inputs: " & " ptr_deref_281_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_281_root_address) & " ptr_deref_281_word_offset_1 = "& Convert_SLV_To_Hex_String(ptr_deref_281_word_offset_1));
          --
        end if; 
        if ptr_deref_281_addr_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_addr_1:finished:  outputs: " & " ptr_deref_281_word_address_1= "  & Convert_SLV_To_Hex_String(ptr_deref_281_word_address_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (33) : ptr_deref_281_addr_1 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_281_root_address;
      ptr_deref_281_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_281_addr_1_req_0;
      ptr_deref_281_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_281_addr_1_req_1;
      ptr_deref_281_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- logger for split-operator ptr_deref_281_addr_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_281_addr_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_addr_2:started:   inputs: " & " ptr_deref_281_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_281_root_address) & " ptr_deref_281_word_offset_2 = "& Convert_SLV_To_Hex_String(ptr_deref_281_word_offset_2));
          --
        end if; 
        if ptr_deref_281_addr_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_addr_2:finished:  outputs: " & " ptr_deref_281_word_address_2= "  & Convert_SLV_To_Hex_String(ptr_deref_281_word_address_2));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (34) : ptr_deref_281_addr_2 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_281_root_address;
      ptr_deref_281_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_281_addr_2_req_0;
      ptr_deref_281_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_281_addr_2_req_1;
      ptr_deref_281_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- logger for split-operator ptr_deref_281_addr_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_281_addr_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_addr_3:started:   inputs: " & " ptr_deref_281_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_281_root_address) & " ptr_deref_281_word_offset_3 = "& Convert_SLV_To_Hex_String(ptr_deref_281_word_offset_3));
          --
        end if; 
        if ptr_deref_281_addr_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_addr_3:finished:  outputs: " & " ptr_deref_281_word_address_3= "  & Convert_SLV_To_Hex_String(ptr_deref_281_word_address_3));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (35) : ptr_deref_281_addr_3 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_281_root_address;
      ptr_deref_281_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_281_addr_3_req_0;
      ptr_deref_281_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_281_addr_3_req_1;
      ptr_deref_281_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- logger for split-operator ptr_deref_87_addr_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_87_addr_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_addr_0:started:   inputs: " & " ptr_deref_87_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_87_root_address) & " ptr_deref_87_word_offset_0 = "& Convert_SLV_To_Hex_String(ptr_deref_87_word_offset_0));
          --
        end if; 
        if ptr_deref_87_addr_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_addr_0:finished:  outputs: " & " ptr_deref_87_word_address_0= "  & Convert_SLV_To_Hex_String(ptr_deref_87_word_address_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (36) : ptr_deref_87_addr_0 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_87_root_address;
      ptr_deref_87_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_87_addr_0_req_0;
      ptr_deref_87_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_87_addr_0_req_1;
      ptr_deref_87_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- logger for split-operator ptr_deref_87_addr_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_87_addr_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_addr_1:started:   inputs: " & " ptr_deref_87_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_87_root_address) & " ptr_deref_87_word_offset_1 = "& Convert_SLV_To_Hex_String(ptr_deref_87_word_offset_1));
          --
        end if; 
        if ptr_deref_87_addr_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_addr_1:finished:  outputs: " & " ptr_deref_87_word_address_1= "  & Convert_SLV_To_Hex_String(ptr_deref_87_word_address_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (37) : ptr_deref_87_addr_1 
    ApIntAdd_group_37: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_87_root_address;
      ptr_deref_87_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_87_addr_1_req_0;
      ptr_deref_87_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_87_addr_1_req_1;
      ptr_deref_87_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_37_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_37_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- logger for split-operator ptr_deref_87_addr_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_87_addr_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_addr_2:started:   inputs: " & " ptr_deref_87_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_87_root_address) & " ptr_deref_87_word_offset_2 = "& Convert_SLV_To_Hex_String(ptr_deref_87_word_offset_2));
          --
        end if; 
        if ptr_deref_87_addr_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_addr_2:finished:  outputs: " & " ptr_deref_87_word_address_2= "  & Convert_SLV_To_Hex_String(ptr_deref_87_word_address_2));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (38) : ptr_deref_87_addr_2 
    ApIntAdd_group_38: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_87_root_address;
      ptr_deref_87_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_87_addr_2_req_0;
      ptr_deref_87_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_87_addr_2_req_1;
      ptr_deref_87_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_38_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_38_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- logger for split-operator ptr_deref_87_addr_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_87_addr_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_addr_3:started:   inputs: " & " ptr_deref_87_root_address = "& Convert_SLV_To_Hex_String(ptr_deref_87_root_address) & " ptr_deref_87_word_offset_3 = "& Convert_SLV_To_Hex_String(ptr_deref_87_word_offset_3));
          --
        end if; 
        if ptr_deref_87_addr_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_addr_3:finished:  outputs: " & " ptr_deref_87_word_address_3= "  & Convert_SLV_To_Hex_String(ptr_deref_87_word_address_3));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (39) : ptr_deref_87_addr_3 
    ApIntAdd_group_39: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_87_root_address;
      ptr_deref_87_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_87_addr_3_req_0;
      ptr_deref_87_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_87_addr_3_req_1;
      ptr_deref_87_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_39_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_39_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_39",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- logger for split-operator type_cast_340_inst flow-through 
    process(type_cast_340_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:type_cast_340_inst:flowthrough inputs: " & " tmp2_336 = "& Convert_SLV_To_Hex_String(tmp2_336) & " outputs:" & " type_cast_340_wire= "  & Convert_SLV_To_Hex_String(type_cast_340_wire));
      --
    end process; 
    -- unary operator type_cast_340_inst
    process(tmp2_336) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp2_336, tmp_var);
      type_cast_340_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator ptr_deref_281_load_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_281_load_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_load_2:started:   inputs: " & " ptr_deref_281_word_address_2 = "& Convert_SLV_To_Hex_String(ptr_deref_281_word_address_2));
          --
        end if; 
        if ptr_deref_281_load_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_load_2:finished:  outputs: " & " ptr_deref_281_data_2= "  & Convert_SLV_To_Hex_String(ptr_deref_281_data_2));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_281_load_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_281_load_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_load_1:started:   inputs: " & " ptr_deref_281_word_address_1 = "& Convert_SLV_To_Hex_String(ptr_deref_281_word_address_1));
          --
        end if; 
        if ptr_deref_281_load_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_load_1:finished:  outputs: " & " ptr_deref_281_data_1= "  & Convert_SLV_To_Hex_String(ptr_deref_281_data_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_212_load_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_212_load_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_load_3:started:   inputs: " & " ptr_deref_212_word_address_3 = "& Convert_SLV_To_Hex_String(ptr_deref_212_word_address_3));
          --
        end if; 
        if ptr_deref_212_load_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_load_3:finished:  outputs: " & " ptr_deref_212_data_3= "  & Convert_SLV_To_Hex_String(ptr_deref_212_data_3));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_281_load_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_281_load_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_load_3:started:   inputs: " & " ptr_deref_281_word_address_3 = "& Convert_SLV_To_Hex_String(ptr_deref_281_word_address_3));
          --
        end if; 
        if ptr_deref_281_load_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_load_3:finished:  outputs: " & " ptr_deref_281_data_3= "  & Convert_SLV_To_Hex_String(ptr_deref_281_data_3));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_281_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_281_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_load_0:started:   inputs: " & " ptr_deref_281_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_281_word_address_0));
          --
        end if; 
        if ptr_deref_281_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_281_load_0:finished:  outputs: " & " ptr_deref_281_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_281_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_212_load_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_212_load_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_load_2:started:   inputs: " & " ptr_deref_212_word_address_2 = "& Convert_SLV_To_Hex_String(ptr_deref_212_word_address_2));
          --
        end if; 
        if ptr_deref_212_load_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_load_2:finished:  outputs: " & " ptr_deref_212_data_2= "  & Convert_SLV_To_Hex_String(ptr_deref_212_data_2));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_212_load_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_212_load_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_load_1:started:   inputs: " & " ptr_deref_212_word_address_1 = "& Convert_SLV_To_Hex_String(ptr_deref_212_word_address_1));
          --
        end if; 
        if ptr_deref_212_load_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_load_1:finished:  outputs: " & " ptr_deref_212_data_1= "  & Convert_SLV_To_Hex_String(ptr_deref_212_data_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_212_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_212_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_load_0:started:   inputs: " & " ptr_deref_212_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_212_word_address_0));
          --
        end if; 
        if ptr_deref_212_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_212_load_0:finished:  outputs: " & " ptr_deref_212_data_0= "  & Convert_SLV_To_Hex_String(ptr_deref_212_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : ptr_deref_281_load_2 ptr_deref_281_load_1 ptr_deref_212_load_3 ptr_deref_281_load_3 ptr_deref_281_load_0 ptr_deref_212_load_2 ptr_deref_212_load_1 ptr_deref_212_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_281_load_2_req_0,
        ptr_deref_281_load_2_ack_0,
        ptr_deref_281_load_2_req_1,
        ptr_deref_281_load_2_ack_1,
        "ptr_deref_281_load_2",
        "memory_space_4" ,
        ptr_deref_281_data_2,
        ptr_deref_281_word_address_2,
        "ptr_deref_281_data_2",
        "ptr_deref_281_word_address_2" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_281_load_1_req_0,
        ptr_deref_281_load_1_ack_0,
        ptr_deref_281_load_1_req_1,
        ptr_deref_281_load_1_ack_1,
        "ptr_deref_281_load_1",
        "memory_space_4" ,
        ptr_deref_281_data_1,
        ptr_deref_281_word_address_1,
        "ptr_deref_281_data_1",
        "ptr_deref_281_word_address_1" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_212_load_3_req_0,
        ptr_deref_212_load_3_ack_0,
        ptr_deref_212_load_3_req_1,
        ptr_deref_212_load_3_ack_1,
        "ptr_deref_212_load_3",
        "memory_space_4" ,
        ptr_deref_212_data_3,
        ptr_deref_212_word_address_3,
        "ptr_deref_212_data_3",
        "ptr_deref_212_word_address_3" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_281_load_3_req_0,
        ptr_deref_281_load_3_ack_0,
        ptr_deref_281_load_3_req_1,
        ptr_deref_281_load_3_ack_1,
        "ptr_deref_281_load_3",
        "memory_space_4" ,
        ptr_deref_281_data_3,
        ptr_deref_281_word_address_3,
        "ptr_deref_281_data_3",
        "ptr_deref_281_word_address_3" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_281_load_0_req_0,
        ptr_deref_281_load_0_ack_0,
        ptr_deref_281_load_0_req_1,
        ptr_deref_281_load_0_ack_1,
        "ptr_deref_281_load_0",
        "memory_space_4" ,
        ptr_deref_281_data_0,
        ptr_deref_281_word_address_0,
        "ptr_deref_281_data_0",
        "ptr_deref_281_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_212_load_2_req_0,
        ptr_deref_212_load_2_ack_0,
        ptr_deref_212_load_2_req_1,
        ptr_deref_212_load_2_ack_1,
        "ptr_deref_212_load_2",
        "memory_space_4" ,
        ptr_deref_212_data_2,
        ptr_deref_212_word_address_2,
        "ptr_deref_212_data_2",
        "ptr_deref_212_word_address_2" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_212_load_1_req_0,
        ptr_deref_212_load_1_ack_0,
        ptr_deref_212_load_1_req_1,
        ptr_deref_212_load_1_ack_1,
        "ptr_deref_212_load_1",
        "memory_space_4" ,
        ptr_deref_212_data_1,
        ptr_deref_212_word_address_1,
        "ptr_deref_212_data_1",
        "ptr_deref_212_word_address_1" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_212_load_0_req_0,
        ptr_deref_212_load_0_ack_0,
        ptr_deref_212_load_0_req_1,
        ptr_deref_212_load_0_ack_1,
        "ptr_deref_212_load_0",
        "memory_space_4" ,
        ptr_deref_212_data_0,
        ptr_deref_212_word_address_0,
        "ptr_deref_212_data_0",
        "ptr_deref_212_word_address_0" -- 
      );
      reqL_unguarded(7) <= ptr_deref_281_load_2_req_0;
      reqL_unguarded(6) <= ptr_deref_281_load_1_req_0;
      reqL_unguarded(5) <= ptr_deref_212_load_3_req_0;
      reqL_unguarded(4) <= ptr_deref_281_load_3_req_0;
      reqL_unguarded(3) <= ptr_deref_281_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_212_load_2_req_0;
      reqL_unguarded(1) <= ptr_deref_212_load_1_req_0;
      reqL_unguarded(0) <= ptr_deref_212_load_0_req_0;
      ptr_deref_281_load_2_ack_0 <= ackL_unguarded(7);
      ptr_deref_281_load_1_ack_0 <= ackL_unguarded(6);
      ptr_deref_212_load_3_ack_0 <= ackL_unguarded(5);
      ptr_deref_281_load_3_ack_0 <= ackL_unguarded(4);
      ptr_deref_281_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_212_load_2_ack_0 <= ackL_unguarded(2);
      ptr_deref_212_load_1_ack_0 <= ackL_unguarded(1);
      ptr_deref_212_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_281_load_2_req_1;
      reqR_unguarded(6) <= ptr_deref_281_load_1_req_1;
      reqR_unguarded(5) <= ptr_deref_212_load_3_req_1;
      reqR_unguarded(4) <= ptr_deref_281_load_3_req_1;
      reqR_unguarded(3) <= ptr_deref_281_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_212_load_2_req_1;
      reqR_unguarded(1) <= ptr_deref_212_load_1_req_1;
      reqR_unguarded(0) <= ptr_deref_212_load_0_req_1;
      ptr_deref_281_load_2_ack_1 <= ackR_unguarded(7);
      ptr_deref_281_load_1_ack_1 <= ackR_unguarded(6);
      ptr_deref_212_load_3_ack_1 <= ackR_unguarded(5);
      ptr_deref_281_load_3_ack_1 <= ackR_unguarded(4);
      ptr_deref_281_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_212_load_2_ack_1 <= ackR_unguarded(2);
      ptr_deref_212_load_1_ack_1 <= ackR_unguarded(1);
      ptr_deref_212_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_281_word_address_2 & ptr_deref_281_word_address_1 & ptr_deref_212_word_address_3 & ptr_deref_281_word_address_3 & ptr_deref_281_word_address_0 & ptr_deref_212_word_address_2 & ptr_deref_212_word_address_1 & ptr_deref_212_word_address_0;
      ptr_deref_281_data_2 <= data_out(63 downto 56);
      ptr_deref_281_data_1 <= data_out(55 downto 48);
      ptr_deref_212_data_3 <= data_out(47 downto 40);
      ptr_deref_281_data_3 <= data_out(39 downto 32);
      ptr_deref_281_data_0 <= data_out(31 downto 24);
      ptr_deref_212_data_2 <= data_out(23 downto 16);
      ptr_deref_212_data_1 <= data_out(15 downto 8);
      ptr_deref_212_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 9,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(8 downto 0),
          mtag => memory_space_4_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(7 downto 0),
          mtag => memory_space_4_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator ptr_deref_184_store_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_184_store_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_store_3:started:   inputs: " & " ptr_deref_184_word_address_3 = "& Convert_SLV_To_Hex_String(ptr_deref_184_word_address_3) & " ptr_deref_184_data_3 = "& Convert_SLV_To_Hex_String(ptr_deref_184_data_3));
          --
        end if; 
        if ptr_deref_184_store_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_store_3:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_184_store_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_184_store_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_store_2:started:   inputs: " & " ptr_deref_184_word_address_2 = "& Convert_SLV_To_Hex_String(ptr_deref_184_word_address_2) & " ptr_deref_184_data_2 = "& Convert_SLV_To_Hex_String(ptr_deref_184_data_2));
          --
        end if; 
        if ptr_deref_184_store_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_store_2:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_184_store_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_184_store_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_store_1:started:   inputs: " & " ptr_deref_184_word_address_1 = "& Convert_SLV_To_Hex_String(ptr_deref_184_word_address_1) & " ptr_deref_184_data_1 = "& Convert_SLV_To_Hex_String(ptr_deref_184_data_1));
          --
        end if; 
        if ptr_deref_184_store_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_store_1:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_184_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_184_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_store_0:started:   inputs: " & " ptr_deref_184_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_184_word_address_0) & " ptr_deref_184_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_184_data_0));
          --
        end if; 
        if ptr_deref_184_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_184_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_87_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_87_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_store_0:started:   inputs: " & " ptr_deref_87_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_87_word_address_0) & " ptr_deref_87_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_87_data_0));
          --
        end if; 
        if ptr_deref_87_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_87_store_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_87_store_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_store_1:started:   inputs: " & " ptr_deref_87_word_address_1 = "& Convert_SLV_To_Hex_String(ptr_deref_87_word_address_1) & " ptr_deref_87_data_1 = "& Convert_SLV_To_Hex_String(ptr_deref_87_data_1));
          --
        end if; 
        if ptr_deref_87_store_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_store_1:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_87_store_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_87_store_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_store_2:started:   inputs: " & " ptr_deref_87_word_address_2 = "& Convert_SLV_To_Hex_String(ptr_deref_87_word_address_2) & " ptr_deref_87_data_2 = "& Convert_SLV_To_Hex_String(ptr_deref_87_data_2));
          --
        end if; 
        if ptr_deref_87_store_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_store_2:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_87_store_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_87_store_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_store_3:started:   inputs: " & " ptr_deref_87_word_address_3 = "& Convert_SLV_To_Hex_String(ptr_deref_87_word_address_3) & " ptr_deref_87_data_3 = "& Convert_SLV_To_Hex_String(ptr_deref_87_data_3));
          --
        end if; 
        if ptr_deref_87_store_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_87_store_3:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_98_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_98_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_98_store_0:started:   inputs: " & " ptr_deref_98_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_98_word_address_0) & " ptr_deref_98_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_98_data_0));
          --
        end if; 
        if ptr_deref_98_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_98_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_109_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_109_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_store_0:started:   inputs: " & " ptr_deref_109_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_109_word_address_0) & " ptr_deref_109_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_109_data_0));
          --
        end if; 
        if ptr_deref_109_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_109_store_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_109_store_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_store_1:started:   inputs: " & " ptr_deref_109_word_address_1 = "& Convert_SLV_To_Hex_String(ptr_deref_109_word_address_1) & " ptr_deref_109_data_1 = "& Convert_SLV_To_Hex_String(ptr_deref_109_data_1));
          --
        end if; 
        if ptr_deref_109_store_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_store_1:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_109_store_2
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_109_store_2_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_store_2:started:   inputs: " & " ptr_deref_109_word_address_2 = "& Convert_SLV_To_Hex_String(ptr_deref_109_word_address_2) & " ptr_deref_109_data_2 = "& Convert_SLV_To_Hex_String(ptr_deref_109_data_2));
          --
        end if; 
        if ptr_deref_109_store_2_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_store_2:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_109_store_3
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_109_store_3_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_store_3:started:   inputs: " & " ptr_deref_109_word_address_3 = "& Convert_SLV_To_Hex_String(ptr_deref_109_word_address_3) & " ptr_deref_109_data_3 = "& Convert_SLV_To_Hex_String(ptr_deref_109_data_3));
          --
        end if; 
        if ptr_deref_109_store_3_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_109_store_3:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_184_store_3_req_0,
      ptr_deref_184_store_3_ack_0,
      ptr_deref_184_store_3_req_1,
      ptr_deref_184_store_3_ack_1,
      "ptr_deref_184_store_3",
      "memory_space_4" ,
      ptr_deref_184_data_3,
      ptr_deref_184_word_address_3,
      "ptr_deref_184_data_3",
      "ptr_deref_184_word_address_3" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_184_store_2_req_0,
      ptr_deref_184_store_2_ack_0,
      ptr_deref_184_store_2_req_1,
      ptr_deref_184_store_2_ack_1,
      "ptr_deref_184_store_2",
      "memory_space_4" ,
      ptr_deref_184_data_2,
      ptr_deref_184_word_address_2,
      "ptr_deref_184_data_2",
      "ptr_deref_184_word_address_2" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_184_store_1_req_0,
      ptr_deref_184_store_1_ack_0,
      ptr_deref_184_store_1_req_1,
      ptr_deref_184_store_1_ack_1,
      "ptr_deref_184_store_1",
      "memory_space_4" ,
      ptr_deref_184_data_1,
      ptr_deref_184_word_address_1,
      "ptr_deref_184_data_1",
      "ptr_deref_184_word_address_1" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_184_store_0_req_0,
      ptr_deref_184_store_0_ack_0,
      ptr_deref_184_store_0_req_1,
      ptr_deref_184_store_0_ack_1,
      "ptr_deref_184_store_0",
      "memory_space_4" ,
      ptr_deref_184_data_0,
      ptr_deref_184_word_address_0,
      "ptr_deref_184_data_0",
      "ptr_deref_184_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_87_store_0_req_0,
      ptr_deref_87_store_0_ack_0,
      ptr_deref_87_store_0_req_1,
      ptr_deref_87_store_0_ack_1,
      "ptr_deref_87_store_0",
      "memory_space_4" ,
      ptr_deref_87_data_0,
      ptr_deref_87_word_address_0,
      "ptr_deref_87_data_0",
      "ptr_deref_87_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_87_store_1_req_0,
      ptr_deref_87_store_1_ack_0,
      ptr_deref_87_store_1_req_1,
      ptr_deref_87_store_1_ack_1,
      "ptr_deref_87_store_1",
      "memory_space_4" ,
      ptr_deref_87_data_1,
      ptr_deref_87_word_address_1,
      "ptr_deref_87_data_1",
      "ptr_deref_87_word_address_1" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_87_store_2_req_0,
      ptr_deref_87_store_2_ack_0,
      ptr_deref_87_store_2_req_1,
      ptr_deref_87_store_2_ack_1,
      "ptr_deref_87_store_2",
      "memory_space_4" ,
      ptr_deref_87_data_2,
      ptr_deref_87_word_address_2,
      "ptr_deref_87_data_2",
      "ptr_deref_87_word_address_2" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_87_store_3_req_0,
      ptr_deref_87_store_3_ack_0,
      ptr_deref_87_store_3_req_1,
      ptr_deref_87_store_3_ack_1,
      "ptr_deref_87_store_3",
      "memory_space_4" ,
      ptr_deref_87_data_3,
      ptr_deref_87_word_address_3,
      "ptr_deref_87_data_3",
      "ptr_deref_87_word_address_3" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_98_store_0_req_0,
      ptr_deref_98_store_0_ack_0,
      ptr_deref_98_store_0_req_1,
      ptr_deref_98_store_0_ack_1,
      "ptr_deref_98_store_0",
      "memory_space_4" ,
      ptr_deref_98_data_0,
      ptr_deref_98_word_address_0,
      "ptr_deref_98_data_0",
      "ptr_deref_98_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_109_store_0_req_0,
      ptr_deref_109_store_0_ack_0,
      ptr_deref_109_store_0_req_1,
      ptr_deref_109_store_0_ack_1,
      "ptr_deref_109_store_0",
      "memory_space_4" ,
      ptr_deref_109_data_0,
      ptr_deref_109_word_address_0,
      "ptr_deref_109_data_0",
      "ptr_deref_109_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_109_store_1_req_0,
      ptr_deref_109_store_1_ack_0,
      ptr_deref_109_store_1_req_1,
      ptr_deref_109_store_1_ack_1,
      "ptr_deref_109_store_1",
      "memory_space_4" ,
      ptr_deref_109_data_1,
      ptr_deref_109_word_address_1,
      "ptr_deref_109_data_1",
      "ptr_deref_109_word_address_1" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_109_store_2_req_0,
      ptr_deref_109_store_2_ack_0,
      ptr_deref_109_store_2_req_1,
      ptr_deref_109_store_2_ack_1,
      "ptr_deref_109_store_2",
      "memory_space_4" ,
      ptr_deref_109_data_2,
      ptr_deref_109_word_address_2,
      "ptr_deref_109_data_2",
      "ptr_deref_109_word_address_2" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_109_store_3_req_0,
      ptr_deref_109_store_3_ack_0,
      ptr_deref_109_store_3_req_1,
      ptr_deref_109_store_3_ack_1,
      "ptr_deref_109_store_3",
      "memory_space_4" ,
      ptr_deref_109_data_3,
      ptr_deref_109_word_address_3,
      "ptr_deref_109_data_3",
      "ptr_deref_109_word_address_3" -- 
    );
    -- shared store operator group (0) : ptr_deref_184_store_3 ptr_deref_184_store_2 ptr_deref_184_store_1 ptr_deref_184_store_0 ptr_deref_87_store_0 ptr_deref_87_store_1 ptr_deref_87_store_2 ptr_deref_87_store_3 ptr_deref_98_store_0 ptr_deref_109_store_0 ptr_deref_109_store_1 ptr_deref_109_store_2 ptr_deref_109_store_3 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(116 downto 0);
      signal data_in: std_logic_vector(103 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 12 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 12 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 12 downto 0);
      signal guard_vector : std_logic_vector( 12 downto 0);
      constant inBUFs : IntegerArray(12 downto 0) := (12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(12 downto 0) := (12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(12 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false);
      constant guardBuffering: IntegerArray(12 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2);
      -- 
    begin -- 
      reqL_unguarded(12) <= ptr_deref_184_store_3_req_0;
      reqL_unguarded(11) <= ptr_deref_184_store_2_req_0;
      reqL_unguarded(10) <= ptr_deref_184_store_1_req_0;
      reqL_unguarded(9) <= ptr_deref_184_store_0_req_0;
      reqL_unguarded(8) <= ptr_deref_87_store_0_req_0;
      reqL_unguarded(7) <= ptr_deref_87_store_1_req_0;
      reqL_unguarded(6) <= ptr_deref_87_store_2_req_0;
      reqL_unguarded(5) <= ptr_deref_87_store_3_req_0;
      reqL_unguarded(4) <= ptr_deref_98_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_109_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_109_store_1_req_0;
      reqL_unguarded(1) <= ptr_deref_109_store_2_req_0;
      reqL_unguarded(0) <= ptr_deref_109_store_3_req_0;
      ptr_deref_184_store_3_ack_0 <= ackL_unguarded(12);
      ptr_deref_184_store_2_ack_0 <= ackL_unguarded(11);
      ptr_deref_184_store_1_ack_0 <= ackL_unguarded(10);
      ptr_deref_184_store_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_87_store_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_87_store_1_ack_0 <= ackL_unguarded(7);
      ptr_deref_87_store_2_ack_0 <= ackL_unguarded(6);
      ptr_deref_87_store_3_ack_0 <= ackL_unguarded(5);
      ptr_deref_98_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_109_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_109_store_1_ack_0 <= ackL_unguarded(2);
      ptr_deref_109_store_2_ack_0 <= ackL_unguarded(1);
      ptr_deref_109_store_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(12) <= ptr_deref_184_store_3_req_1;
      reqR_unguarded(11) <= ptr_deref_184_store_2_req_1;
      reqR_unguarded(10) <= ptr_deref_184_store_1_req_1;
      reqR_unguarded(9) <= ptr_deref_184_store_0_req_1;
      reqR_unguarded(8) <= ptr_deref_87_store_0_req_1;
      reqR_unguarded(7) <= ptr_deref_87_store_1_req_1;
      reqR_unguarded(6) <= ptr_deref_87_store_2_req_1;
      reqR_unguarded(5) <= ptr_deref_87_store_3_req_1;
      reqR_unguarded(4) <= ptr_deref_98_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_109_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_109_store_1_req_1;
      reqR_unguarded(1) <= ptr_deref_109_store_2_req_1;
      reqR_unguarded(0) <= ptr_deref_109_store_3_req_1;
      ptr_deref_184_store_3_ack_1 <= ackR_unguarded(12);
      ptr_deref_184_store_2_ack_1 <= ackR_unguarded(11);
      ptr_deref_184_store_1_ack_1 <= ackR_unguarded(10);
      ptr_deref_184_store_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_87_store_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_87_store_1_ack_1 <= ackR_unguarded(7);
      ptr_deref_87_store_2_ack_1 <= ackR_unguarded(6);
      ptr_deref_87_store_3_ack_1 <= ackR_unguarded(5);
      ptr_deref_98_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_109_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_109_store_1_ack_1 <= ackR_unguarded(2);
      ptr_deref_109_store_2_ack_1 <= ackR_unguarded(1);
      ptr_deref_109_store_3_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_6: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_7: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_8: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_9: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_10: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_11: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_12: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 13, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_184_word_address_3 & ptr_deref_184_word_address_2 & ptr_deref_184_word_address_1 & ptr_deref_184_word_address_0 & ptr_deref_87_word_address_0 & ptr_deref_87_word_address_1 & ptr_deref_87_word_address_2 & ptr_deref_87_word_address_3 & ptr_deref_98_word_address_0 & ptr_deref_109_word_address_0 & ptr_deref_109_word_address_1 & ptr_deref_109_word_address_2 & ptr_deref_109_word_address_3;
      data_in <= ptr_deref_184_data_3 & ptr_deref_184_data_2 & ptr_deref_184_data_1 & ptr_deref_184_data_0 & ptr_deref_87_data_0 & ptr_deref_87_data_1 & ptr_deref_87_data_2 & ptr_deref_87_data_3 & ptr_deref_98_data_0 & ptr_deref_109_data_0 & ptr_deref_109_data_1 & ptr_deref_109_data_2 & ptr_deref_109_data_3;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 9,
        data_width => 8,
        num_reqs => 13,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(8 downto 0),
          mdata => memory_space_4_sr_data(7 downto 0),
          mtag => memory_space_4_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 13,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logger for split-operator ptr_deref_195_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_195_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_195_store_0:started:   inputs: " & " ptr_deref_195_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_195_word_address_0) & " ptr_deref_195_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_195_data_0));
          --
        end if; 
        if ptr_deref_195_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_195_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator ptr_deref_120_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ptr_deref_120_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_120_store_0:started:   inputs: " & " ptr_deref_120_word_address_0 = "& Convert_SLV_To_Hex_String(ptr_deref_120_word_address_0) & " ptr_deref_120_data_0 = "& Convert_SLV_To_Hex_String(ptr_deref_120_data_0));
          --
        end if; 
        if ptr_deref_120_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:ptr_deref_120_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_195_store_0_req_0,
      ptr_deref_195_store_0_ack_0,
      ptr_deref_195_store_0_req_1,
      ptr_deref_195_store_0_ack_1,
      "ptr_deref_195_store_0",
      "memory_space_3" ,
      ptr_deref_195_data_0,
      ptr_deref_195_word_address_0,
      "ptr_deref_195_data_0",
      "ptr_deref_195_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_120_store_0_req_0,
      ptr_deref_120_store_0_ack_0,
      ptr_deref_120_store_0_req_1,
      ptr_deref_120_store_0_ack_1,
      "ptr_deref_120_store_0",
      "memory_space_3" ,
      ptr_deref_120_data_0,
      ptr_deref_120_word_address_0,
      "ptr_deref_120_data_0",
      "ptr_deref_120_word_address_0" -- 
    );
    -- shared store operator group (1) : ptr_deref_195_store_0 ptr_deref_120_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_195_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_120_store_0_req_0;
      ptr_deref_195_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_120_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_195_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_120_store_0_req_1;
      ptr_deref_195_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_120_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_195_word_address_0 & ptr_deref_120_word_address_0;
      data_in <= ptr_deref_195_data_0 & ptr_deref_120_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(6 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- logger for split-operator RPIPE_maxpool_input_pipe_188_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_188_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:RPIPE_maxpool_input_pipe_188_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_188_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:RPIPE_maxpool_input_pipe_188_inst:finished:  outputs: " & " call3_189= "  & Convert_SLV_To_Hex_String(call3_189));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator RPIPE_maxpool_input_pipe_177_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_maxpool_input_pipe_177_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:RPIPE_maxpool_input_pipe_177_inst:started:   PipeRead from maxpool_input_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_maxpool_input_pipe_177_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:RPIPE_maxpool_input_pipe_177_inst:finished:  outputs: " & " call_178= "  & Convert_SLV_To_Hex_String(call_178));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_188_inst RPIPE_maxpool_input_pipe_177_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_188_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_177_inst_req_0;
      RPIPE_maxpool_input_pipe_188_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_177_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_188_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_177_inst_req_1;
      RPIPE_maxpool_input_pipe_188_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_177_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      call3_189 <= data_out(31 downto 16);
      call_178 <= data_out(15 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 16,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator call_stmt_373_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_373_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:call_stmt_373_call:started:  Call to module fill_T inputs: " & " iNsTr_22_364 = "& Convert_SLV_To_Hex_String(iNsTr_22_364));
          --
        end if; 
        if call_stmt_373_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:testConfigure:DP:call_stmt_373_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_373_call 
    fill_T_call_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_373_call_req_0;
      call_stmt_373_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_373_call_req_1;
      call_stmt_373_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      fill_T_call_group_0_gI: SplitGuardInterface generic map(name => "fill_T_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_22_364;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => fill_T_call_reqs(0),
          ackR => fill_T_call_acks(0),
          dataR => fill_T_call_data(63 downto 0),
          tagR => fill_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => fill_T_return_acks(0), -- cross-over
          ackL => fill_T_return_reqs(0), -- cross-over
          tagL => fill_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_1802_start: Boolean;
  signal timer_CP_1802_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_401_load_0_req_1 : boolean;
  signal LOAD_count_401_load_0_ack_1 : boolean;
  signal LOAD_count_401_load_0_ack_0 : boolean;
  signal LOAD_count_401_load_0_req_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_1802_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1802_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_1802_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1802_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,timer_CP_1802_start,"timer cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,timer_CP_1802_symbol, "timer cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_1802: Block -- control-path 
    signal timer_CP_1802_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_1802_elements(0) <= timer_CP_1802_start;
    timer_CP_1802_symbol <= timer_CP_1802_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_update_start_
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_sample_start_
      -- CP-element group 0: 	 assign_stmt_402/$entry
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_Update/$entry
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_402/LOAD_count_401_Update/word_access_complete/$entry
      -- 
    -- logger for CP element group timer_CP_1802_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timer_CP_1802_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:timer_CP_1802_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:LOAD_count_401_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:LOAD_count_401_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1802_elements(0), ack => LOAD_count_401_load_0_req_0); -- 
    cr_1834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1802_elements(0), ack => LOAD_count_401_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_402/LOAD_count_401_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_402/LOAD_count_401_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_402/LOAD_count_401_sample_completed_
      -- CP-element group 1: 	 assign_stmt_402/LOAD_count_401_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_402/LOAD_count_401_Sample/word_access_start/word_0/$exit
      -- 
    -- logger for CP element group timer_CP_1802_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timer_CP_1802_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:timer_CP_1802_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:LOAD_count_401_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_401_load_0_ack_0, ack => timer_CP_1802_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_402/LOAD_count_401_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_402/LOAD_count_401_Update/LOAD_count_401_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_402/LOAD_count_401_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_402/LOAD_count_401_update_completed_
      -- CP-element group 2: 	 assign_stmt_402/LOAD_count_401_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_402/$exit
      -- CP-element group 2: 	 assign_stmt_402/LOAD_count_401_Update/LOAD_count_401_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_402/LOAD_count_401_Update/LOAD_count_401_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_402/LOAD_count_401_Update/$exit
      -- CP-element group 2: 	 assign_stmt_402/LOAD_count_401_Update/LOAD_count_401_Merge/merge_ack
      -- 
    -- logger for CP element group timer_CP_1802_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timer_CP_1802_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:timer_CP_1802_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timer:CP:LOAD_count_401_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_401_load_0_ack_1, ack => timer_CP_1802_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_401_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_401_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_401_word_address_0 <= "0";
    -- logger for operator LOAD_count_401_gather_scatter flow-through 
    process(c_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:timer:DP:LOAD_count_401_gather_scatter:flowthrough  inputs: " & " LOAD_count_401_data_0 = "& Convert_SLV_To_Hex_String(LOAD_count_401_data_0) & "outputs: " & " c_buffer= "  & Convert_SLV_To_Hex_String(c_buffer));
      --
    end process; 
    -- equivalence LOAD_count_401_gather_scatter
    process(LOAD_count_401_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_401_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- logger for split-operator LOAD_count_401_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_count_401_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timer:DP:LOAD_count_401_load_0:started:   inputs: " & " LOAD_count_401_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_count_401_word_address_0));
          --
        end if; 
        if LOAD_count_401_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timer:DP:LOAD_count_401_load_0:finished:  outputs: " & " LOAD_count_401_data_0= "  & Convert_SLV_To_Hex_String(LOAD_count_401_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : LOAD_count_401_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_count_401_load_0_req_0,
        LOAD_count_401_load_0_ack_0,
        LOAD_count_401_load_0_req_1,
        LOAD_count_401_load_0_ack_1,
        "LOAD_count_401_load_0",
        "memory_space_2" ,
        LOAD_count_401_data_0,
        LOAD_count_401_word_address_0,
        "LOAD_count_401_data_0",
        "LOAD_count_401_word_address_0" -- 
      );
      reqL_unguarded(0) <= LOAD_count_401_load_0_req_0;
      LOAD_count_401_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_401_load_0_req_1;
      LOAD_count_401_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_401_word_address_0;
      LOAD_count_401_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_5245_start: Boolean;
  signal timerDaemon_CP_5245_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal STORE_count_2067_store_0_req_0 : boolean;
  signal STORE_count_2067_store_0_ack_0 : boolean;
  signal ADD_u64_u64_2065_inst_req_0 : boolean;
  signal ADD_u64_u64_2065_inst_ack_0 : boolean;
  signal ADD_u64_u64_2065_inst_req_1 : boolean;
  signal ADD_u64_u64_2065_inst_ack_1 : boolean;
  signal STORE_count_2067_store_0_req_1 : boolean;
  signal do_while_stmt_2057_branch_req_0 : boolean;
  signal phi_stmt_2059_req_1 : boolean;
  signal phi_stmt_2059_req_0 : boolean;
  signal phi_stmt_2059_ack_0 : boolean;
  signal STORE_count_2067_store_0_ack_1 : boolean;
  signal do_while_stmt_2057_branch_ack_0 : boolean;
  signal do_while_stmt_2057_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_5245_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_5245_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_5245_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_5245_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,timerDaemon_CP_5245_start,"timerDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,timerDaemon_CP_5245_symbol, "timerDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_5245: Block -- control-path 
    signal timerDaemon_CP_5245_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_5245_elements(0) <= timerDaemon_CP_5245_start;
    timerDaemon_CP_5245_symbol <= timerDaemon_CP_5245_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2056/$entry
      -- CP-element group 0: 	 branch_block_stmt_2056/branch_block_stmt_2056__entry__
      -- CP-element group 0: 	 branch_block_stmt_2056/do_while_stmt_2057__entry__
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2056/$exit
      -- CP-element group 1: 	 branch_block_stmt_2056/branch_block_stmt_2056__exit__
      -- CP-element group 1: 	 branch_block_stmt_2056/do_while_stmt_2057__exit__
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_5245_elements(1) <= timerDaemon_CP_5245_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2056/do_while_stmt_2057/$entry
      -- CP-element group 2: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057__entry__
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_5245_elements(2) <= timerDaemon_CP_5245_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057__exit__
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2056/do_while_stmt_2057/loop_back
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2056/do_while_stmt_2057/condition_done
      -- CP-element group 5: 	 branch_block_stmt_2056/do_while_stmt_2057/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_2056/do_while_stmt_2057/loop_taken/$entry
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_5245_elements(5) <= timerDaemon_CP_5245_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2056/do_while_stmt_2057/loop_body_done
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_5245_elements(6) <= timerDaemon_CP_5245_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_5245_elements(7) <= timerDaemon_CP_5245_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_5245_elements(8) <= timerDaemon_CP_5245_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	35 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/loop_body_start
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	35 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/condition_evaluated
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:do_while_stmt_2057_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_5269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_5269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5245_elements(10), ack => do_while_stmt_2057_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5245_elements(15) & timerDaemon_CP_5245_elements(35);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5245_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_sample_start__ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5245_elements(12) & timerDaemon_CP_5245_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5245_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_sample_start_
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5245_elements(9) & timerDaemon_CP_5245_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5245_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_update_start_
      -- CP-element group 13: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_update_start__ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5245_elements(9) & timerDaemon_CP_5245_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5245_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_sample_completed__ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	31 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_update_completed__ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_loopback_trigger
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_5245_elements(16) <= timerDaemon_CP_5245_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_loopback_sample_req_ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:phi_stmt_2059_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_2059_loopback_sample_req_5284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2059_loopback_sample_req_5284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5245_elements(17), ack => phi_stmt_2059_req_1); -- 
    -- Element group timerDaemon_CP_5245_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_entry_trigger
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_5245_elements(18) <= timerDaemon_CP_5245_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_entry_sample_req_ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:phi_stmt_2059_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_2059_entry_sample_req_5287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2059_entry_sample_req_5287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5245_elements(19), ack => phi_stmt_2059_req_0); -- 
    -- Element group timerDaemon_CP_5245_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/phi_stmt_2059_phi_mux_ack_ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:phi_stmt_2059_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_2059_phi_mux_ack_5290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2059_ack_0, ack => timerDaemon_CP_5245_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/type_cast_2062_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/type_cast_2062_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/type_cast_2062_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/type_cast_2062_sample_completed_
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/type_cast_2062_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/type_cast_2062_update_start_
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/type_cast_2062_update_completed__ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_5245_elements(23) <= timerDaemon_CP_5245_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/type_cast_2062_update_completed_
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_5245_elements(22), ack => timerDaemon_CP_5245_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_sample_start__ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_update_start__ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(26) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_Sample/$entry
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:ADD_u64_u64_2065_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5245_elements(27), ack => ADD_u64_u64_2065_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5245_elements(25) & timerDaemon_CP_5245_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5245_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_Update/cr
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:ADD_u64_u64_2065_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_5316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5245_elements(28), ack => ADD_u64_u64_2065_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5245_elements(26) & timerDaemon_CP_5245_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5245_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_sample_completed__ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:ADD_u64_u64_2065_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2065_inst_ack_0, ack => timerDaemon_CP_5245_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/ADD_u64_u64_2065_update_completed__ps
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:ADD_u64_u64_2065_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2065_inst_ack_1, ack => timerDaemon_CP_5245_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/word_access_start/word_0/rr
      -- CP-element group 31: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/STORE_count_2067_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/STORE_count_2067_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/STORE_count_2067_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/STORE_count_2067_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/word_access_start/word_0/$entry
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:STORE_count_2067_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5245_elements(31), ack => STORE_count_2067_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_5245_elements(9) & timerDaemon_CP_5245_elements(15) & timerDaemon_CP_5245_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5245_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Update/word_access_complete/word_0/cr
      -- CP-element group 32: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_update_start_
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:STORE_count_2067_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_5350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5245_elements(32), ack => STORE_count_2067_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_5245_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5245_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/word_access_start/word_0/ra
      -- CP-element group 33: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_sample_completed_
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:STORE_count_2067_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_2067_store_0_ack_0, ack => timerDaemon_CP_5245_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/STORE_count_2067_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:STORE_count_2067_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_2067_store_0_ack_1, ack => timerDaemon_CP_5245_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group timerDaemon_CP_5245_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_5245_elements(9), ack => timerDaemon_CP_5245_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_2056/do_while_stmt_2057/do_while_stmt_2057_loop_body/$exit
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(36) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5245_elements(14) & timerDaemon_CP_5245_elements(34);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5245_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_2056/do_while_stmt_2057/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_2056/do_while_stmt_2057/loop_exit/ack
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:do_while_stmt_2057_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2057_branch_ack_0, ack => timerDaemon_CP_5245_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_2056/do_while_stmt_2057/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_2056/do_while_stmt_2057/loop_taken/ack
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:do_while_stmt_2057_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2057_branch_ack_1, ack => timerDaemon_CP_5245_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_2056/do_while_stmt_2057/$exit
      -- 
    -- logger for CP element group timerDaemon_CP_5245_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and timerDaemon_CP_5245_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:timerDaemon:CP:timerDaemon_CP_5245_elements(39) fired."); 
        -- 
      end if; --
    end process; 
    timerDaemon_CP_5245_elements(39) <= timerDaemon_CP_5245_elements(3);
    timerDaemon_do_while_stmt_2057_terminator_5361: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_2057_terminator_5361", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_5245_elements(6),loop_continue => timerDaemon_CP_5245_elements(38),loop_terminate => timerDaemon_CP_5245_elements(37),loop_back => timerDaemon_CP_5245_elements(4),loop_exit => timerDaemon_CP_5245_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2059_phi_seq_5318_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_5245_elements(18);
      timerDaemon_CP_5245_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_5245_elements(21);
      timerDaemon_CP_5245_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_5245_elements(23);
      timerDaemon_CP_5245_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_5245_elements(16);
      timerDaemon_CP_5245_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_5245_elements(29);
      timerDaemon_CP_5245_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_5245_elements(30);
      timerDaemon_CP_5245_elements(17) <= phi_mux_reqs(1);
      phi_stmt_2059_phi_seq_5318 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_2059_phi_seq_5318") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_5245_elements(11), 
          phi_sample_ack => timerDaemon_CP_5245_elements(14), 
          phi_update_req => timerDaemon_CP_5245_elements(13), 
          phi_update_ack => timerDaemon_CP_5245_elements(15), 
          phi_mux_ack => timerDaemon_CP_5245_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_5270_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_5245_elements(7);
        preds(1)  <= timerDaemon_CP_5245_elements(8);
        entry_tmerge_5270 : transition_merge -- 
          generic map(name => " entry_tmerge_5270")
          port map (preds => preds, symbol_out => timerDaemon_CP_5245_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_2065_wire : std_logic_vector(63 downto 0);
    signal STORE_count_2067_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_2067_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_2064_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2071_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_2059 : std_logic_vector(63 downto 0);
    signal type_cast_2062_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_2067_word_address_0 <= "0";
    konst_2064_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_2071_wire_constant <= "1";
    type_cast_2062_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- logger for phi phi_stmt_2059
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_2059_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:timerDaemon:DP:phi_stmt_2059:input-0 type_cast_2062_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_2062_wire_constant));
          --
        end if;
        if phi_stmt_2059_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:timerDaemon:DP:phi_stmt_2059:input-1 ADD_u64_u64_2065_wire= " & Convert_SLV_To_Hex_String(ADD_u64_u64_2065_wire));
          --
        end if;
        if phi_stmt_2059_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:timerDaemon:DP:phi_stmt_2059:sample-completed");
          --
        end if;
        if phi_stmt_2059_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:timerDaemon:DP:phi_stmt_2059:output ncount_2059= " & Convert_SLV_To_Hex_String(ncount_2059));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_2059: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2062_wire_constant & ADD_u64_u64_2065_wire;
      req <= phi_stmt_2059_req_0 & phi_stmt_2059_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2059",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2059_ack_0,
          idata => idata,
          odata => ncount_2059,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2059
    -- logger for operator STORE_count_2067_gather_scatter flow-through 
    process(STORE_count_2067_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:timerDaemon:DP:STORE_count_2067_gather_scatter:flowthrough  inputs: " & " ncount_2059 = "& Convert_SLV_To_Hex_String(ncount_2059) & "outputs: " & " STORE_count_2067_data_0= "  & Convert_SLV_To_Hex_String(STORE_count_2067_data_0));
      --
    end process; 
    -- equivalence STORE_count_2067_gather_scatter
    process(ncount_2059) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_2059;
      ov(63 downto 0) := iv;
      STORE_count_2067_data_0 <= ov(63 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_2057_branch_req_0," req0 do_while_stmt_2057_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_2057_branch_ack_0," ack0 do_while_stmt_2057_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_2057_branch_ack_1," ack1 do_while_stmt_2057_branch");
    do_while_stmt_2057_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2071_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2057_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2057_branch_req_0,
          ack0 => do_while_stmt_2057_branch_ack_0,
          ack1 => do_while_stmt_2057_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u64_u64_2065_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u64_u64_2065_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timerDaemon:DP:ADD_u64_u64_2065_inst:started:   inputs: " & " ncount_2059 = "& Convert_SLV_To_Hex_String(ncount_2059) & " konst_2064_wire_constant = "& Convert_SLV_To_Hex_String(konst_2064_wire_constant));
          --
        end if; 
        if ADD_u64_u64_2065_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timerDaemon:DP:ADD_u64_u64_2065_inst:finished:  outputs: " & " ADD_u64_u64_2065_wire= "  & Convert_SLV_To_Hex_String(ADD_u64_u64_2065_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : ADD_u64_u64_2065_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_2059;
      ADD_u64_u64_2065_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2065_inst_req_0;
      ADD_u64_u64_2065_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2065_inst_req_1;
      ADD_u64_u64_2065_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator STORE_count_2067_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_count_2067_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timerDaemon:DP:STORE_count_2067_store_0:started:   inputs: " & " STORE_count_2067_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_count_2067_word_address_0) & " STORE_count_2067_data_0 = "& Convert_SLV_To_Hex_String(STORE_count_2067_data_0));
          --
        end if; 
        if STORE_count_2067_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:timerDaemon:DP:STORE_count_2067_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_count_2067_store_0_req_0,
      STORE_count_2067_store_0_ack_0,
      STORE_count_2067_store_0_req_1,
      STORE_count_2067_store_0_ack_1,
      "STORE_count_2067_store_0",
      "memory_space_2" ,
      STORE_count_2067_data_0,
      STORE_count_2067_word_address_0,
      "STORE_count_2067_data_0",
      "STORE_count_2067_word_address_0" -- 
    );
    -- shared store operator group (0) : STORE_count_2067_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_2067_store_0_req_0;
      STORE_count_2067_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_2067_store_0_req_1;
      STORE_count_2067_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_2067_word_address_0;
      data_in <= STORE_count_2067_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(15 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(15 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(255 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(37 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(17 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(41 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(8 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module fill_T
  component fill_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module fill_T
  signal fill_T_addr :  std_logic_vector(63 downto 0);
  signal fill_T_in_args    : std_logic_vector(63 downto 0);
  signal fill_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal fill_T_tag_out   : std_logic_vector(1 downto 0);
  signal fill_T_start_req : std_logic;
  signal fill_T_start_ack : std_logic;
  signal fill_T_fin_req   : std_logic;
  signal fill_T_fin_ack : std_logic;
  -- caller side aggregated signals for module fill_T
  signal fill_T_call_reqs: std_logic_vector(0 downto 0);
  signal fill_T_call_acks: std_logic_vector(0 downto 0);
  signal fill_T_return_reqs: std_logic_vector(0 downto 0);
  signal fill_T_return_acks: std_logic_vector(0 downto 0);
  signal fill_T_call_data: std_logic_vector(63 downto 0);
  signal fill_T_call_tag: std_logic_vector(0 downto 0);
  signal fill_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module maxPool3D
  component maxPool3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_call_acks : in   std_logic_vector(0 downto 0);
      maxPool4_call_data : out  std_logic_vector(159 downto 0);
      maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
      maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_return_acks : in   std_logic_vector(0 downto 0);
      maxPool4_return_data : in   std_logic_vector(7 downto 0);
      maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
      sendB_call_reqs : out  std_logic_vector(0 downto 0);
      sendB_call_acks : in   std_logic_vector(0 downto 0);
      sendB_call_tag  :  out  std_logic_vector(0 downto 0);
      sendB_return_reqs : out  std_logic_vector(0 downto 0);
      sendB_return_acks : in   std_logic_vector(0 downto 0);
      sendB_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool3D
  signal maxPool3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool3D_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool3D_start_req : std_logic;
  signal maxPool3D_start_ack : std_logic;
  signal maxPool3D_fin_req   : std_logic;
  signal maxPool3D_fin_ack : std_logic;
  -- declarations related to module maxPool4
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      output : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool4
  signal maxPool4_addr :  std_logic_vector(31 downto 0);
  signal maxPool4_addr1 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr2 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr3 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr4 :  std_logic_vector(31 downto 0);
  signal maxPool4_output :  std_logic_vector(7 downto 0);
  signal maxPool4_in_args    : std_logic_vector(159 downto 0);
  signal maxPool4_out_args   : std_logic_vector(7 downto 0);
  signal maxPool4_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool4_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool4_start_req : std_logic;
  signal maxPool4_start_ack : std_logic;
  signal maxPool4_fin_req   : std_logic;
  signal maxPool4_fin_ack : std_logic;
  -- caller side aggregated signals for module maxPool4
  signal maxPool4_call_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_call_acks: std_logic_vector(0 downto 0);
  signal maxPool4_return_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_return_acks: std_logic_vector(0 downto 0);
  signal maxPool4_call_data: std_logic_vector(159 downto 0);
  signal maxPool4_call_tag: std_logic_vector(0 downto 0);
  signal maxPool4_return_data: std_logic_vector(7 downto 0);
  signal maxPool4_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendB
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendB
  signal sendB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendB_tag_out   : std_logic_vector(1 downto 0);
  signal sendB_start_req : std_logic;
  signal sendB_start_ack : std_logic;
  signal sendB_fin_req   : std_logic;
  signal sendB_fin_ack : std_logic;
  -- caller side aggregated signals for module sendB
  signal sendB_call_reqs: std_logic_vector(0 downto 0);
  signal sendB_call_acks: std_logic_vector(0 downto 0);
  signal sendB_return_reqs: std_logic_vector(0 downto 0);
  signal sendB_return_acks: std_logic_vector(0 downto 0);
  signal sendB_call_tag: std_logic_vector(0 downto 0);
  signal sendB_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(8 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      fill_T_call_reqs : out  std_logic_vector(0 downto 0);
      fill_T_call_acks : in   std_logic_vector(0 downto 0);
      fill_T_call_data : out  std_logic_vector(63 downto 0);
      fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
      fill_T_return_reqs : out  std_logic_vector(0 downto 0);
      fill_T_return_acks : in   std_logic_vector(0 downto 0);
      fill_T_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module fill_T
  fill_T_addr <= fill_T_in_args(63 downto 0);
  -- call arbiter for module fill_T
  fill_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => fill_T_call_reqs,
      call_acks => fill_T_call_acks,
      return_reqs => fill_T_return_reqs,
      return_acks => fill_T_return_acks,
      call_data  => fill_T_call_data,
      call_tag  => fill_T_call_tag,
      return_tag  => fill_T_return_tag,
      call_mtag => fill_T_tag_in,
      return_mtag => fill_T_tag_out,
      call_mreq => fill_T_start_req,
      call_mack => fill_T_start_ack,
      return_mreq => fill_T_fin_req,
      return_mack => fill_T_fin_ack,
      call_mdata => fill_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  fill_T_instance:fill_T-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => fill_T_addr,
      start_req => fill_T_start_req,
      start_ack => fill_T_start_ack,
      fin_req => fill_T_fin_req,
      fin_ack => fill_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(255 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(19 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(1 downto 1),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(1 downto 1),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(31 downto 16),
      tag_in => fill_T_tag_in,
      tag_out => fill_T_tag_out-- 
    ); -- 
  -- module maxPool3D
  maxPool3D_instance:maxPool3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => maxPool3D_start_req,
      start_ack => maxPool3D_start_ack,
      fin_req => maxPool3D_fin_req,
      fin_ack => maxPool3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(6 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(1 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(8 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(20 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(7 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(3 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      maxPool4_call_reqs => maxPool4_call_reqs(0 downto 0),
      maxPool4_call_acks => maxPool4_call_acks(0 downto 0),
      maxPool4_call_data => maxPool4_call_data(159 downto 0),
      maxPool4_call_tag => maxPool4_call_tag(0 downto 0),
      maxPool4_return_reqs => maxPool4_return_reqs(0 downto 0),
      maxPool4_return_acks => maxPool4_return_acks(0 downto 0),
      maxPool4_return_data => maxPool4_return_data(7 downto 0),
      maxPool4_return_tag => maxPool4_return_tag(0 downto 0),
      sendB_call_reqs => sendB_call_reqs(0 downto 0),
      sendB_call_acks => sendB_call_acks(0 downto 0),
      sendB_call_tag => sendB_call_tag(0 downto 0),
      sendB_return_reqs => sendB_return_reqs(0 downto 0),
      sendB_return_acks => sendB_return_acks(0 downto 0),
      sendB_return_tag => sendB_return_tag(0 downto 0),
      tag_in => maxPool3D_tag_in,
      tag_out => maxPool3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  maxPool3D_tag_in <= (others => '0');
  maxPool3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => maxPool3D_start_req, start_ack => maxPool3D_start_ack,  fin_req => maxPool3D_fin_req,  fin_ack => maxPool3D_fin_ack);
  -- module maxPool4
  maxPool4_addr <= maxPool4_in_args(159 downto 128);
  maxPool4_addr1 <= maxPool4_in_args(127 downto 96);
  maxPool4_addr2 <= maxPool4_in_args(95 downto 64);
  maxPool4_addr3 <= maxPool4_in_args(63 downto 32);
  maxPool4_addr4 <= maxPool4_in_args(31 downto 0);
  maxPool4_out_args <= maxPool4_output ;
  -- call arbiter for module maxPool4
  maxPool4_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 160,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => maxPool4_call_reqs,
      call_acks => maxPool4_call_acks,
      return_reqs => maxPool4_return_reqs,
      return_acks => maxPool4_return_acks,
      call_data  => maxPool4_call_data,
      call_tag  => maxPool4_call_tag,
      return_tag  => maxPool4_return_tag,
      call_mtag => maxPool4_tag_in,
      return_mtag => maxPool4_tag_out,
      return_data =>maxPool4_return_data,
      call_mreq => maxPool4_start_req,
      call_mack => maxPool4_start_ack,
      return_mreq => maxPool4_fin_req,
      return_mack => maxPool4_fin_ack,
      call_mdata => maxPool4_in_args,
      return_mdata => maxPool4_out_args,
      clk => clk, 
      reset => reset --
    ); --
  maxPool4_instance:maxPool4-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => maxPool4_addr,
      addr1 => maxPool4_addr1,
      addr2 => maxPool4_addr2,
      addr3 => maxPool4_addr3,
      addr4 => maxPool4_addr4,
      output => maxPool4_output,
      start_req => maxPool4_start_req,
      start_ack => maxPool4_start_ack,
      fin_req => maxPool4_fin_req,
      fin_ack => maxPool4_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(19 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      tag_in => maxPool4_tag_in,
      tag_out => maxPool4_tag_out-- 
    ); -- 
  -- module sendB
  -- call arbiter for module sendB
  sendB_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendB_call_reqs,
      call_acks => sendB_call_acks,
      return_reqs => sendB_return_reqs,
      return_acks => sendB_return_acks,
      call_tag  => sendB_call_tag,
      return_tag  => sendB_return_tag,
      call_mtag => sendB_tag_in,
      return_mtag => sendB_tag_out,
      call_mreq => sendB_start_req,
      call_mack => sendB_start_ack,
      return_mreq => sendB_fin_req,
      return_mack => sendB_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendB_instance:sendB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendB_start_req,
      start_ack => sendB_start_ack,
      fin_req => sendB_fin_req,
      fin_ack => sendB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 7),
      memory_space_3_lr_tag => memory_space_3_lr_tag(37 downto 19),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 32),
      memory_space_3_lc_tag => memory_space_3_lc_tag(3 downto 2),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 0),
      tag_in => sendB_tag_in,
      tag_out => sendB_tag_out-- 
    ); -- 
  -- module testConfigure
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_4_lr_req => memory_space_4_lr_req(1 downto 1),
      memory_space_4_lr_ack => memory_space_4_lr_ack(1 downto 1),
      memory_space_4_lr_addr => memory_space_4_lr_addr(17 downto 9),
      memory_space_4_lr_tag => memory_space_4_lr_tag(41 downto 21),
      memory_space_4_lc_req => memory_space_4_lc_req(1 downto 1),
      memory_space_4_lc_ack => memory_space_4_lc_ack(1 downto 1),
      memory_space_4_lc_data => memory_space_4_lc_data(15 downto 8),
      memory_space_4_lc_tag => memory_space_4_lc_tag(7 downto 4),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(6 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(31 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(8 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(7 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(20 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(3 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(15 downto 0),
      fill_T_call_reqs => fill_T_call_reqs(0 downto 0),
      fill_T_call_acks => fill_T_call_acks(0 downto 0),
      fill_T_call_data => fill_T_call_data(63 downto 0),
      fill_T_call_tag => fill_T_call_tag(0 downto 0),
      fill_T_return_reqs => fill_T_return_reqs(0 downto 0),
      fill_T_return_acks => fill_T_return_acks(0 downto 0),
      fill_T_return_tag => fill_T_return_tag(0 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 2,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 256,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 256
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 2,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 2,
      num_stores => 1,
      addr_width => 9,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 9,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
