-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_3910_start: Boolean;
  signal convTranspose_CP_3910_symbol: Boolean;
  -- volatile/operator module components. 
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_Block0_done_1347_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1337_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1356_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1347_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1334_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1334_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1356_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1334_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1343_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1356_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1343_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1353_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1337_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1353_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1356_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1343_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1343_inst_req_0 : boolean;
  signal call_stmt_1332_call_ack_1 : boolean;
  signal call_stmt_1332_call_req_1 : boolean;
  signal call_stmt_1332_call_ack_0 : boolean;
  signal call_stmt_1332_call_req_0 : boolean;
  signal RPIPE_Block1_done_1350_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1350_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1340_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1340_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1350_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1340_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1350_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1340_inst_req_0 : boolean;
  signal call_stmt_1359_call_ack_1 : boolean;
  signal call_stmt_1359_call_req_1 : boolean;
  signal call_stmt_1359_call_ack_0 : boolean;
  signal call_stmt_1359_call_req_0 : boolean;
  signal WPIPE_Block1_start_1337_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1337_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1334_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1347_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1353_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1347_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1353_inst_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_3910_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3910_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_3910_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3910_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_3910: Block -- control-path 
    signal convTranspose_CP_3910_elements: BooleanArray(21 downto 0);
    -- 
  begin -- 
    convTranspose_CP_3910_elements(0) <= convTranspose_CP_3910_start;
    convTranspose_CP_3910_symbol <= convTranspose_CP_3910_elements(21);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_1330/branch_block_stmt_1330__entry__
      -- CP-element group 0: 	 branch_block_stmt_1330/call_stmt_1332/$entry
      -- CP-element group 0: 	 branch_block_stmt_1330/$entry
      -- CP-element group 0: 	 branch_block_stmt_1330/call_stmt_1332__entry__
      -- CP-element group 0: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_Update/ccr
      -- CP-element group 0: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_sample_start_
      -- CP-element group 0: 	 $entry
      -- 
    ccr_3941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(0), ack => call_stmt_1332_call_req_1); -- 
    crr_3936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(0), ack => call_stmt_1332_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_sample_completed_
      -- 
    cra_3937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1332_call_ack_0, ack => convTranspose_CP_3910_elements(1)); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (31) 
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357__entry__
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1330/call_stmt_1332__exit__
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/$entry
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1330/call_stmt_1332/call_stmt_1332_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1330/call_stmt_1332/$exit
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_sample_start_
      -- 
    cca_3942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1332_call_ack_1, ack => convTranspose_CP_3910_elements(2)); -- 
    rr_4009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => RPIPE_Block0_done_1347_inst_req_0); -- 
    req_3953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => WPIPE_Block0_start_1334_inst_req_0); -- 
    rr_4051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => RPIPE_Block3_done_1356_inst_req_0); -- 
    rr_4037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => RPIPE_Block2_done_1353_inst_req_0); -- 
    req_3995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => WPIPE_Block3_start_1343_inst_req_0); -- 
    rr_4023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => RPIPE_Block1_done_1350_inst_req_0); -- 
    req_3981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => WPIPE_Block2_start_1340_inst_req_0); -- 
    req_3967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => WPIPE_Block1_start_1337_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_Update/req
      -- CP-element group 3: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_Sample/ack
      -- 
    ack_3954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1334_inst_ack_0, ack => convTranspose_CP_3910_elements(3)); -- 
    req_3958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(3), ack => WPIPE_Block0_start_1334_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	19 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_Update/ack
      -- CP-element group 4: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block0_start_1334_update_completed_
      -- 
    ack_3959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1334_inst_ack_1, ack => convTranspose_CP_3910_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_Update/req
      -- CP-element group 5: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_Sample/ack
      -- CP-element group 5: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_Sample/$exit
      -- 
    ack_3968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1337_inst_ack_0, ack => convTranspose_CP_3910_elements(5)); -- 
    req_3972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(5), ack => WPIPE_Block1_start_1337_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	19 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block1_start_1337_update_completed_
      -- 
    ack_3973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1337_inst_ack_1, ack => convTranspose_CP_3910_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_Update/req
      -- CP-element group 7: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_Sample/ack
      -- CP-element group 7: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_sample_completed_
      -- 
    ack_3982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1340_inst_ack_0, ack => convTranspose_CP_3910_elements(7)); -- 
    req_3986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(7), ack => WPIPE_Block2_start_1340_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	19 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_Update/ack
      -- CP-element group 8: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block2_start_1340_update_completed_
      -- 
    ack_3987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1340_inst_ack_1, ack => convTranspose_CP_3910_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_Update/req
      -- CP-element group 9: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_Sample/ack
      -- CP-element group 9: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_sample_completed_
      -- 
    ack_3996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1343_inst_ack_0, ack => convTranspose_CP_3910_elements(9)); -- 
    req_4000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(9), ack => WPIPE_Block3_start_1343_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	19 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_Update/ack
      -- CP-element group 10: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/WPIPE_Block3_start_1343_update_completed_
      -- 
    ack_4001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1343_inst_ack_1, ack => convTranspose_CP_3910_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_Update/$entry
      -- 
    ra_4010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1347_inst_ack_0, ack => convTranspose_CP_3910_elements(11)); -- 
    cr_4014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(11), ack => RPIPE_Block0_done_1347_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	19 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block0_done_1347_Update/$exit
      -- 
    ca_4015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1347_inst_ack_1, ack => convTranspose_CP_3910_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_Sample/$exit
      -- 
    ra_4024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1350_inst_ack_0, ack => convTranspose_CP_3910_elements(13)); -- 
    cr_4028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(13), ack => RPIPE_Block1_done_1350_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	19 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block1_done_1350_Update/$exit
      -- 
    ca_4029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1350_inst_ack_1, ack => convTranspose_CP_3910_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_Update/cr
      -- 
    ra_4038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1353_inst_ack_0, ack => convTranspose_CP_3910_elements(15)); -- 
    cr_4042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(15), ack => RPIPE_Block2_done_1353_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	19 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block2_done_1353_Update/ca
      -- 
    ca_4043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1353_inst_ack_1, ack => convTranspose_CP_3910_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_update_start_
      -- 
    ra_4052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1356_inst_ack_0, ack => convTranspose_CP_3910_elements(17)); -- 
    cr_4056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(17), ack => RPIPE_Block3_done_1356_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/RPIPE_Block3_done_1356_update_completed_
      -- 
    ca_4057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1356_inst_ack_1, ack => convTranspose_CP_3910_elements(18)); -- 
    -- CP-element group 19:  join  fork  transition  place  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	8 
    -- CP-element group 19: 	10 
    -- CP-element group 19: 	12 
    -- CP-element group 19: 	6 
    -- CP-element group 19: 	4 
    -- CP-element group 19: 	18 
    -- CP-element group 19: 	14 
    -- CP-element group 19: 	16 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (10) 
      -- CP-element group 19: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357__exit__
      -- CP-element group 19: 	 branch_block_stmt_1330/call_stmt_1359__entry__
      -- CP-element group 19: 	 branch_block_stmt_1330/assign_stmt_1336_to_assign_stmt_1357/$exit
      -- CP-element group 19: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1330/call_stmt_1359/$entry
      -- CP-element group 19: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_Update/ccr
      -- CP-element group 19: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_Sample/crr
      -- 
    ccr_4073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(19), ack => call_stmt_1359_call_req_1); -- 
    crr_4068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(19), ack => call_stmt_1359_call_req_0); -- 
    convTranspose_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= convTranspose_CP_3910_elements(8) & convTranspose_CP_3910_elements(10) & convTranspose_CP_3910_elements(12) & convTranspose_CP_3910_elements(6) & convTranspose_CP_3910_elements(4) & convTranspose_CP_3910_elements(18) & convTranspose_CP_3910_elements(14) & convTranspose_CP_3910_elements(16);
      gj_convTranspose_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3910_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_Sample/cra
      -- CP-element group 20: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_Sample/$exit
      -- 
    cra_4069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1359_call_ack_0, ack => convTranspose_CP_3910_elements(20)); -- 
    -- CP-element group 21:  transition  place  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (16) 
      -- CP-element group 21: 	 branch_block_stmt_1330/branch_block_stmt_1330__exit__
      -- CP-element group 21: 	 branch_block_stmt_1330/merge_stmt_1361_PhiAck/dummy
      -- CP-element group 21: 	 branch_block_stmt_1330/merge_stmt_1361_PhiReqMerge
      -- CP-element group 21: 	 branch_block_stmt_1330/merge_stmt_1361__exit__
      -- CP-element group 21: 	 branch_block_stmt_1330/return__
      -- CP-element group 21: 	 branch_block_stmt_1330/call_stmt_1359__exit__
      -- CP-element group 21: 	 branch_block_stmt_1330/merge_stmt_1361_PhiAck/$exit
      -- CP-element group 21: 	 branch_block_stmt_1330/$exit
      -- CP-element group 21: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1330/return___PhiReq/$exit
      -- CP-element group 21: 	 branch_block_stmt_1330/return___PhiReq/$entry
      -- CP-element group 21: 	 branch_block_stmt_1330/call_stmt_1359/$exit
      -- CP-element group 21: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_Update/cca
      -- CP-element group 21: 	 branch_block_stmt_1330/call_stmt_1359/call_stmt_1359_Update/$exit
      -- CP-element group 21: 	 $exit
      -- CP-element group 21: 	 branch_block_stmt_1330/merge_stmt_1361_PhiAck/$entry
      -- 
    cca_4074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1359_call_ack_1, ack => convTranspose_CP_3910_elements(21)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call11_1357 : std_logic_vector(15 downto 0);
    signal call5_1348 : std_logic_vector(15 downto 0);
    signal call7_1351 : std_logic_vector(15 downto 0);
    signal call9_1354 : std_logic_vector(15 downto 0);
    signal call_1332 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    -- shared inport operator group (0) : RPIPE_Block0_done_1347_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1347_inst_req_0;
      RPIPE_Block0_done_1347_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1347_inst_req_1;
      RPIPE_Block0_done_1347_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call5_1348 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1350_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1350_inst_req_0;
      RPIPE_Block1_done_1350_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1350_inst_req_1;
      RPIPE_Block1_done_1350_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call7_1351 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1353_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1353_inst_req_0;
      RPIPE_Block2_done_1353_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1353_inst_req_1;
      RPIPE_Block2_done_1353_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call9_1354 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1356_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1356_inst_req_0;
      RPIPE_Block3_done_1356_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1356_inst_req_1;
      RPIPE_Block3_done_1356_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call11_1357 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_Block0_start_1334_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_start_1334_inst_req_0;
      WPIPE_Block0_start_1334_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_start_1334_inst_req_1;
      WPIPE_Block0_start_1334_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1332;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1337_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_start_1337_inst_req_0;
      WPIPE_Block1_start_1337_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_start_1337_inst_req_1;
      WPIPE_Block1_start_1337_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1332;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1340_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_start_1340_inst_req_0;
      WPIPE_Block2_start_1340_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_start_1340_inst_req_1;
      WPIPE_Block2_start_1340_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1332;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1343_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_start_1343_inst_req_0;
      WPIPE_Block3_start_1343_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_start_1343_inst_req_1;
      WPIPE_Block3_start_1343_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1332;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_stmt_1332_call 
    testConfigure_call_group_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1332_call_req_0;
      call_stmt_1332_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1332_call_req_1;
      call_stmt_1332_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_1332 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1359_call 
    sendOutput_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1359_call_req_0;
      call_stmt_1359_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1359_call_req_1;
      call_stmt_1359_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_4083_start: Boolean;
  signal convTransposeA_CP_4083_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1680_inst_ack_0 : boolean;
  signal array_obj_ref_1717_index_offset_req_0 : boolean;
  signal ptr_deref_1475_load_0_ack_1 : boolean;
  signal addr_of_1687_final_reg_req_1 : boolean;
  signal type_cast_1680_inst_ack_1 : boolean;
  signal ptr_deref_1691_load_0_ack_0 : boolean;
  signal ptr_deref_1691_load_0_req_1 : boolean;
  signal type_cast_1680_inst_req_1 : boolean;
  signal ptr_deref_1493_load_0_ack_0 : boolean;
  signal type_cast_1680_inst_req_0 : boolean;
  signal addr_of_1687_final_reg_ack_1 : boolean;
  signal array_obj_ref_1717_index_offset_ack_0 : boolean;
  signal ptr_deref_1691_load_0_ack_1 : boolean;
  signal ptr_deref_1493_load_0_req_0 : boolean;
  signal type_cast_1711_inst_ack_0 : boolean;
  signal type_cast_1711_inst_req_1 : boolean;
  signal type_cast_1711_inst_ack_1 : boolean;
  signal ptr_deref_1691_load_0_req_0 : boolean;
  signal type_cast_1711_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1367_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1367_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1367_inst_req_1 : boolean;
  signal array_obj_ref_1686_index_offset_ack_1 : boolean;
  signal RPIPE_Block0_start_1367_inst_ack_1 : boolean;
  signal ptr_deref_1475_load_0_req_1 : boolean;
  signal array_obj_ref_1686_index_offset_req_1 : boolean;
  signal type_cast_1649_inst_ack_1 : boolean;
  signal type_cast_1649_inst_req_1 : boolean;
  signal array_obj_ref_1686_index_offset_ack_0 : boolean;
  signal type_cast_1649_inst_ack_0 : boolean;
  signal type_cast_1649_inst_req_0 : boolean;
  signal ptr_deref_1380_load_0_req_0 : boolean;
  signal ptr_deref_1380_load_0_ack_0 : boolean;
  signal ptr_deref_1493_load_0_ack_1 : boolean;
  signal ptr_deref_1380_load_0_req_1 : boolean;
  signal ptr_deref_1380_load_0_ack_1 : boolean;
  signal array_obj_ref_1686_index_offset_req_0 : boolean;
  signal addr_of_1687_final_reg_ack_0 : boolean;
  signal type_cast_1527_inst_ack_1 : boolean;
  signal type_cast_1527_inst_req_1 : boolean;
  signal type_cast_1527_inst_ack_0 : boolean;
  signal type_cast_1527_inst_req_0 : boolean;
  signal ptr_deref_1493_load_0_req_1 : boolean;
  signal ptr_deref_1392_load_0_req_0 : boolean;
  signal ptr_deref_1392_load_0_ack_0 : boolean;
  signal ptr_deref_1392_load_0_req_1 : boolean;
  signal ptr_deref_1392_load_0_ack_1 : boolean;
  signal addr_of_1687_final_reg_req_0 : boolean;
  signal type_cast_1522_inst_ack_1 : boolean;
  signal type_cast_1522_inst_req_1 : boolean;
  signal type_cast_1522_inst_ack_0 : boolean;
  signal type_cast_1522_inst_req_0 : boolean;
  signal ptr_deref_1402_load_0_req_0 : boolean;
  signal ptr_deref_1402_load_0_ack_0 : boolean;
  signal ptr_deref_1402_load_0_req_1 : boolean;
  signal ptr_deref_1402_load_0_ack_1 : boolean;
  signal type_cast_1406_inst_req_0 : boolean;
  signal type_cast_1406_inst_ack_0 : boolean;
  signal type_cast_1406_inst_req_1 : boolean;
  signal type_cast_1406_inst_ack_1 : boolean;
  signal ptr_deref_1418_load_0_req_0 : boolean;
  signal ptr_deref_1418_load_0_ack_0 : boolean;
  signal ptr_deref_1418_load_0_req_1 : boolean;
  signal ptr_deref_1418_load_0_ack_1 : boolean;
  signal LOAD_padding_1421_load_0_req_0 : boolean;
  signal LOAD_padding_1421_load_0_ack_0 : boolean;
  signal LOAD_padding_1421_load_0_req_1 : boolean;
  signal LOAD_padding_1421_load_0_ack_1 : boolean;
  signal type_cast_1425_inst_req_0 : boolean;
  signal type_cast_1425_inst_ack_0 : boolean;
  signal type_cast_1425_inst_req_1 : boolean;
  signal type_cast_1425_inst_ack_1 : boolean;
  signal ptr_deref_1435_load_0_req_0 : boolean;
  signal ptr_deref_1435_load_0_ack_0 : boolean;
  signal ptr_deref_1435_load_0_req_1 : boolean;
  signal ptr_deref_1435_load_0_ack_1 : boolean;
  signal type_cast_1439_inst_req_0 : boolean;
  signal type_cast_1439_inst_ack_0 : boolean;
  signal type_cast_1439_inst_req_1 : boolean;
  signal type_cast_1439_inst_ack_1 : boolean;
  signal ptr_deref_1451_load_0_req_0 : boolean;
  signal ptr_deref_1451_load_0_ack_0 : boolean;
  signal ptr_deref_1451_load_0_req_1 : boolean;
  signal ptr_deref_1451_load_0_ack_1 : boolean;
  signal ptr_deref_1463_load_0_req_0 : boolean;
  signal ptr_deref_1463_load_0_ack_0 : boolean;
  signal ptr_deref_1463_load_0_req_1 : boolean;
  signal ptr_deref_1463_load_0_ack_1 : boolean;
  signal ptr_deref_1475_load_0_req_0 : boolean;
  signal ptr_deref_1475_load_0_ack_0 : boolean;
  signal array_obj_ref_1717_index_offset_req_1 : boolean;
  signal array_obj_ref_1717_index_offset_ack_1 : boolean;
  signal addr_of_1718_final_reg_req_0 : boolean;
  signal addr_of_1718_final_reg_ack_0 : boolean;
  signal addr_of_1718_final_reg_req_1 : boolean;
  signal addr_of_1718_final_reg_ack_1 : boolean;
  signal ptr_deref_1721_store_0_req_0 : boolean;
  signal ptr_deref_1721_store_0_ack_0 : boolean;
  signal ptr_deref_1721_store_0_req_1 : boolean;
  signal ptr_deref_1721_store_0_ack_1 : boolean;
  signal type_cast_1727_inst_req_0 : boolean;
  signal type_cast_1727_inst_ack_0 : boolean;
  signal type_cast_1727_inst_req_1 : boolean;
  signal type_cast_1727_inst_ack_1 : boolean;
  signal if_stmt_1740_branch_req_0 : boolean;
  signal if_stmt_1740_branch_ack_1 : boolean;
  signal if_stmt_1740_branch_ack_0 : boolean;
  signal type_cast_1764_inst_req_0 : boolean;
  signal type_cast_1764_inst_ack_0 : boolean;
  signal type_cast_1764_inst_req_1 : boolean;
  signal type_cast_1764_inst_ack_1 : boolean;
  signal type_cast_1773_inst_req_0 : boolean;
  signal type_cast_1773_inst_ack_0 : boolean;
  signal type_cast_1773_inst_req_1 : boolean;
  signal type_cast_1773_inst_ack_1 : boolean;
  signal type_cast_1790_inst_req_0 : boolean;
  signal type_cast_1790_inst_ack_0 : boolean;
  signal type_cast_1790_inst_req_1 : boolean;
  signal type_cast_1790_inst_ack_1 : boolean;
  signal if_stmt_1797_branch_req_0 : boolean;
  signal if_stmt_1797_branch_ack_1 : boolean;
  signal if_stmt_1797_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1805_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1805_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1805_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1805_inst_ack_1 : boolean;
  signal phi_stmt_1503_req_0 : boolean;
  signal phi_stmt_1510_req_0 : boolean;
  signal type_cast_1509_inst_req_0 : boolean;
  signal type_cast_1509_inst_ack_0 : boolean;
  signal type_cast_1509_inst_req_1 : boolean;
  signal type_cast_1509_inst_ack_1 : boolean;
  signal phi_stmt_1503_req_1 : boolean;
  signal type_cast_1516_inst_req_0 : boolean;
  signal type_cast_1516_inst_ack_0 : boolean;
  signal type_cast_1516_inst_req_1 : boolean;
  signal type_cast_1516_inst_ack_1 : boolean;
  signal phi_stmt_1510_req_1 : boolean;
  signal phi_stmt_1503_ack_0 : boolean;
  signal phi_stmt_1510_ack_0 : boolean;
  signal type_cast_1639_inst_req_0 : boolean;
  signal type_cast_1639_inst_ack_0 : boolean;
  signal type_cast_1639_inst_req_1 : boolean;
  signal type_cast_1639_inst_ack_1 : boolean;
  signal phi_stmt_1633_req_1 : boolean;
  signal phi_stmt_1633_req_0 : boolean;
  signal phi_stmt_1633_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_4083_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_4083_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_4083_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_4083_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_4083: Block -- control-path 
    signal convTransposeA_CP_4083_elements: BooleanArray(88 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_4083_elements(0) <= convTransposeA_CP_4083_start;
    convTransposeA_CP_4083_symbol <= convTransposeA_CP_4083_elements(68);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1365/$entry
      -- CP-element group 0: 	 branch_block_stmt_1365/branch_block_stmt_1365__entry__
      -- CP-element group 0: 	 branch_block_stmt_1365/assign_stmt_1368__entry__
      -- CP-element group 0: 	 branch_block_stmt_1365/assign_stmt_1368/$entry
      -- CP-element group 0: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_Sample/rr
      -- 
    rr_4131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(0), ack => RPIPE_Block0_start_1367_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_Update/cr
      -- 
    ra_4132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1367_inst_ack_0, ack => convTransposeA_CP_4083_elements(1)); -- 
    cr_4136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(1), ack => RPIPE_Block0_start_1367_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1368__exit__
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500__entry__
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1368/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1368/RPIPE_Block0_start_1367_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Sample/word_access_start/word_0/rr
      -- 
    ca_4137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1367_inst_ack_1, ack => convTransposeA_CP_4083_elements(2)); -- 
    rr_4648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1493_load_0_req_0); -- 
    cr_4609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1475_load_0_req_1); -- 
    rr_4173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1380_load_0_req_0); -- 
    cr_4184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1380_load_0_req_1); -- 
    cr_4659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1493_load_0_req_1); -- 
    rr_4223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1392_load_0_req_0); -- 
    cr_4234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1392_load_0_req_1); -- 
    rr_4273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1402_load_0_req_0); -- 
    cr_4284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1402_load_0_req_1); -- 
    cr_4303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => type_cast_1406_inst_req_1); -- 
    rr_4337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1418_load_0_req_0); -- 
    cr_4348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1418_load_0_req_1); -- 
    rr_4370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => LOAD_padding_1421_load_0_req_0); -- 
    cr_4381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => LOAD_padding_1421_load_0_req_1); -- 
    cr_4400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => type_cast_1425_inst_req_1); -- 
    rr_4434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1435_load_0_req_0); -- 
    cr_4445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1435_load_0_req_1); -- 
    cr_4464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => type_cast_1439_inst_req_1); -- 
    rr_4498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1451_load_0_req_0); -- 
    cr_4509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1451_load_0_req_1); -- 
    rr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1463_load_0_req_0); -- 
    cr_4559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1463_load_0_req_1); -- 
    rr_4598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1475_load_0_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Sample/word_access_start/word_0/ra
      -- 
    ra_4174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1380_load_0_ack_0, ack => convTransposeA_CP_4083_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	29 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/ptr_deref_1380_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/ptr_deref_1380_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/ptr_deref_1380_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1380_Update/ptr_deref_1380_Merge/merge_ack
      -- 
    ca_4185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1380_load_0_ack_1, ack => convTransposeA_CP_4083_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Sample/word_access_start/word_0/ra
      -- 
    ra_4224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1392_load_0_ack_0, ack => convTransposeA_CP_4083_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	29 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/ptr_deref_1392_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/ptr_deref_1392_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/ptr_deref_1392_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1392_Update/ptr_deref_1392_Merge/merge_ack
      -- 
    ca_4235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1392_load_0_ack_1, ack => convTransposeA_CP_4083_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Sample/word_access_start/word_0/ra
      -- 
    ra_4274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1402_load_0_ack_0, ack => convTransposeA_CP_4083_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/ptr_deref_1402_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/ptr_deref_1402_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/ptr_deref_1402_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1402_Update/ptr_deref_1402_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_Sample/rr
      -- 
    ca_4285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1402_load_0_ack_1, ack => convTransposeA_CP_4083_elements(8)); -- 
    rr_4298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(8), ack => type_cast_1406_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_Sample/ra
      -- 
    ra_4299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_0, ack => convTransposeA_CP_4083_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1406_Update/ca
      -- 
    ca_4304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_1, ack => convTransposeA_CP_4083_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Sample/word_access_start/word_0/ra
      -- 
    ra_4338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1418_load_0_ack_0, ack => convTransposeA_CP_4083_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/ptr_deref_1418_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/ptr_deref_1418_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/ptr_deref_1418_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1418_Update/ptr_deref_1418_Merge/merge_ack
      -- 
    ca_4349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1418_load_0_ack_1, ack => convTransposeA_CP_4083_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Sample/word_access_start/word_0/ra
      -- 
    ra_4371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1421_load_0_ack_0, ack => convTransposeA_CP_4083_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/LOAD_padding_1421_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/LOAD_padding_1421_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/LOAD_padding_1421_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/LOAD_padding_1421_Update/LOAD_padding_1421_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_Sample/rr
      -- 
    ca_4382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1421_load_0_ack_1, ack => convTransposeA_CP_4083_elements(14)); -- 
    rr_4395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(14), ack => type_cast_1425_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_Sample/ra
      -- 
    ra_4396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_0, ack => convTransposeA_CP_4083_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1425_Update/ca
      -- 
    ca_4401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_1, ack => convTransposeA_CP_4083_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Sample/word_access_start/word_0/ra
      -- 
    ra_4435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1435_load_0_ack_0, ack => convTransposeA_CP_4083_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (12) 
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/ptr_deref_1435_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/ptr_deref_1435_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/ptr_deref_1435_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1435_Update/ptr_deref_1435_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_Sample/rr
      -- 
    ca_4446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1435_load_0_ack_1, ack => convTransposeA_CP_4083_elements(18)); -- 
    rr_4459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(18), ack => type_cast_1439_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_Sample/ra
      -- 
    ra_4460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1439_inst_ack_0, ack => convTransposeA_CP_4083_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/type_cast_1439_Update/ca
      -- 
    ca_4465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1439_inst_ack_1, ack => convTransposeA_CP_4083_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Sample/word_access_start/word_0/ra
      -- 
    ra_4499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1451_load_0_ack_0, ack => convTransposeA_CP_4083_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/ptr_deref_1451_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/ptr_deref_1451_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/ptr_deref_1451_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1451_Update/ptr_deref_1451_Merge/merge_ack
      -- 
    ca_4510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1451_load_0_ack_1, ack => convTransposeA_CP_4083_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Sample/word_access_start/word_0/ra
      -- 
    ra_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1463_load_0_ack_0, ack => convTransposeA_CP_4083_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/ptr_deref_1463_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/ptr_deref_1463_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/ptr_deref_1463_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1463_Update/ptr_deref_1463_Merge/merge_ack
      -- 
    ca_4560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1463_load_0_ack_1, ack => convTransposeA_CP_4083_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Sample/word_access_start/word_0/ra
      -- 
    ra_4599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1475_load_0_ack_0, ack => convTransposeA_CP_4083_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/ptr_deref_1475_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/ptr_deref_1475_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/ptr_deref_1475_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/ptr_deref_1475_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1475_update_completed_
      -- 
    ca_4610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1475_load_0_ack_1, ack => convTransposeA_CP_4083_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Sample/word_access_start/word_0/ra
      -- CP-element group 27: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Sample/$exit
      -- 
    ra_4649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1493_load_0_ack_0, ack => convTransposeA_CP_4083_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/ptr_deref_1493_Merge/merge_ack
      -- CP-element group 28: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/ptr_deref_1493_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/ptr_deref_1493_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/ptr_deref_1493_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/ptr_deref_1493_Update/word_access_complete/$exit
      -- 
    ca_4660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1493_load_0_ack_1, ack => convTransposeA_CP_4083_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	4 
    -- CP-element group 29: 	6 
    -- CP-element group 29: 	10 
    -- CP-element group 29: 	12 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	69 
    -- CP-element group 29: 	70 
    -- CP-element group 29:  members (8) 
      -- CP-element group 29: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500__exit__
      -- CP-element group 29: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_1365/assign_stmt_1377_to_assign_stmt_1500/$exit
      -- CP-element group 29: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/$entry
      -- CP-element group 29: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/$entry
      -- CP-element group 29: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/$entry
      -- 
    convTransposeA_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(16) & convTransposeA_CP_4083_elements(20) & convTransposeA_CP_4083_elements(22) & convTransposeA_CP_4083_elements(24) & convTransposeA_CP_4083_elements(26) & convTransposeA_CP_4083_elements(28) & convTransposeA_CP_4083_elements(4) & convTransposeA_CP_4083_elements(6) & convTransposeA_CP_4083_elements(10) & convTransposeA_CP_4083_elements(12);
      gj_convTransposeA_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	82 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_Sample/$exit
      -- 
    ra_4677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1522_inst_ack_0, ack => convTransposeA_CP_4083_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	82 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_update_completed_
      -- 
    ca_4682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1522_inst_ack_1, ack => convTransposeA_CP_4083_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	82 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_sample_completed_
      -- 
    ra_4691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1527_inst_ack_0, ack => convTransposeA_CP_4083_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	82 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_update_completed_
      -- 
    ca_4696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1527_inst_ack_1, ack => convTransposeA_CP_4083_elements(33)); -- 
    -- CP-element group 34:  join  transition  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	86 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/$exit
      -- CP-element group 34: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630__exit__
      -- CP-element group 34: 	 branch_block_stmt_1365/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 34: 	 branch_block_stmt_1365/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_1365/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1633/$entry
      -- CP-element group 34: 	 branch_block_stmt_1365/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/$entry
      -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(31) & convTransposeA_CP_4083_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_sample_completed_
      -- 
    ra_4708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1649_inst_ack_0, ack => convTransposeA_CP_4083_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	88 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	45 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_update_completed_
      -- 
    ca_4713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1649_inst_ack_1, ack => convTransposeA_CP_4083_elements(36)); -- 
    rr_4721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(36), ack => type_cast_1680_inst_req_0); -- 
    rr_4831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(36), ack => type_cast_1711_inst_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_sample_completed_
      -- 
    ra_4722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1680_inst_ack_0, ack => convTransposeA_CP_4083_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	88 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (16) 
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_resize_1/$entry
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_resize_1/index_resize_req
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_resize_1/$exit
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_scaled_1
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_computed_1
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_resize_1/index_resize_ack
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_scale_1/$entry
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_resized_1
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_final_index_sum_regn_Sample/req
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_final_index_sum_regn_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_scale_1/scale_rename_ack
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_scale_1/scale_rename_req
      -- CP-element group 38: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_index_scale_1/$exit
      -- 
    ca_4727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1680_inst_ack_1, ack => convTransposeA_CP_4083_elements(38)); -- 
    req_4752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(38), ack => array_obj_ref_1686_index_offset_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	56 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_final_index_sum_regn_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_final_index_sum_regn_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_final_index_sum_regn_sample_complete
      -- 
    ack_4753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1686_index_offset_ack_0, ack => convTransposeA_CP_4083_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	88 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (11) 
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_base_plus_offset/sum_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_request/$entry
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_base_plus_offset/sum_rename_req
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_root_address_calculated
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_offset_calculated
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_base_plus_offset/$exit
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_base_plus_offset/$entry
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_final_index_sum_regn_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_final_index_sum_regn_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_request/req
      -- 
    ack_4758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1686_index_offset_ack_1, ack => convTransposeA_CP_4083_elements(40)); -- 
    req_4767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(40), ack => addr_of_1687_final_reg_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_request/$exit
      -- CP-element group 41: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_request/ack
      -- 
    ack_4768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1687_final_reg_ack_0, ack => convTransposeA_CP_4083_elements(41)); -- 
    -- CP-element group 42:  join  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	88 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (24) 
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_complete/$exit
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_base_addr_resize/$entry
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_base_address_resized
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_complete/ack
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_word_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_base_addr_resize/base_resize_ack
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_word_addrgen/root_register_req
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_word_addrgen/root_register_ack
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Sample/word_access_start/word_0/rr
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Sample/word_access_start/$entry
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_word_addrgen/$exit
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_word_addrgen/$entry
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_base_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_base_addr_resize/base_resize_req
      -- CP-element group 42: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_base_addr_resize/$exit
      -- 
    ack_4773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1687_final_reg_ack_1, ack => convTransposeA_CP_4083_elements(42)); -- 
    rr_4806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(42), ack => ptr_deref_1691_load_0_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Sample/word_access_start/word_0/ra
      -- CP-element group 43: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Sample/word_access_start/$exit
      -- 
    ra_4807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1691_load_0_ack_0, ack => convTransposeA_CP_4083_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	88 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	51 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/ptr_deref_1691_Merge/merge_req
      -- CP-element group 44: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/word_access_complete/word_0/ca
      -- CP-element group 44: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/ptr_deref_1691_Merge/$entry
      -- CP-element group 44: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/ptr_deref_1691_Merge/$exit
      -- CP-element group 44: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/ptr_deref_1691_Merge/merge_ack
      -- CP-element group 44: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_update_completed_
      -- 
    ca_4818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1691_load_0_ack_1, ack => convTransposeA_CP_4083_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	36 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_Sample/$exit
      -- 
    ra_4832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1711_inst_ack_0, ack => convTransposeA_CP_4083_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	88 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (16) 
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_final_index_sum_regn_Sample/req
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_resize_1/index_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_computed_1
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_scale_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_scale_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_resized_1
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_final_index_sum_regn_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_scale_1/scale_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_resize_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_resize_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_resize_1/index_resize_req
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_scaled_1
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_index_scale_1/scale_rename_req
      -- CP-element group 46: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_Update/$exit
      -- 
    ca_4837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1711_inst_ack_1, ack => convTransposeA_CP_4083_elements(46)); -- 
    req_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(46), ack => array_obj_ref_1717_index_offset_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_final_index_sum_regn_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_final_index_sum_regn_Sample/ack
      -- CP-element group 47: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_final_index_sum_regn_sample_complete
      -- 
    ack_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1717_index_offset_ack_0, ack => convTransposeA_CP_4083_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	88 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (11) 
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_offset_calculated
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_final_index_sum_regn_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_request/$entry
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_final_index_sum_regn_Update/ack
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_request/req
      -- 
    ack_4868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1717_index_offset_ack_1, ack => convTransposeA_CP_4083_elements(48)); -- 
    req_4877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(48), ack => addr_of_1718_final_reg_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_request/$exit
      -- CP-element group 49: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_request/ack
      -- 
    ack_4878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1718_final_reg_ack_0, ack => convTransposeA_CP_4083_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	88 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (19) 
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_word_addrgen/root_register_ack
      -- 
    ack_4883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1718_final_reg_ack_1, ack => convTransposeA_CP_4083_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	44 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/ptr_deref_1721_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/ptr_deref_1721_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/ptr_deref_1721_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/ptr_deref_1721_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/word_access_start/word_0/rr
      -- 
    rr_4921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(51), ack => ptr_deref_1721_store_0_req_0); -- 
    convTransposeA_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(44) & convTransposeA_CP_4083_elements(50);
      gj_convTransposeA_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Sample/word_access_start/word_0/ra
      -- 
    ra_4922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1721_store_0_ack_0, ack => convTransposeA_CP_4083_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	88 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Update/word_access_complete/word_0/ca
      -- 
    ca_4933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1721_store_0_ack_1, ack => convTransposeA_CP_4083_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	88 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_Sample/ra
      -- 
    ra_4942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1727_inst_ack_0, ack => convTransposeA_CP_4083_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	88 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_Update/ca
      -- 
    ca_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1727_inst_ack_1, ack => convTransposeA_CP_4083_elements(55)); -- 
    -- CP-element group 56:  branch  join  transition  place  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: 	47 
    -- CP-element group 56: 	53 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (10) 
      -- CP-element group 56: 	 branch_block_stmt_1365/R_cmp_1741_place
      -- CP-element group 56: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739__exit__
      -- CP-element group 56: 	 branch_block_stmt_1365/if_stmt_1740__entry__
      -- CP-element group 56: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/$exit
      -- CP-element group 56: 	 branch_block_stmt_1365/if_stmt_1740_dead_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1365/if_stmt_1740_eval_test/$entry
      -- CP-element group 56: 	 branch_block_stmt_1365/if_stmt_1740_eval_test/$exit
      -- CP-element group 56: 	 branch_block_stmt_1365/if_stmt_1740_eval_test/branch_req
      -- CP-element group 56: 	 branch_block_stmt_1365/if_stmt_1740_if_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1365/if_stmt_1740_else_link/$entry
      -- 
    branch_req_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(56), ack => if_stmt_1740_branch_req_0); -- 
    convTransposeA_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(39) & convTransposeA_CP_4083_elements(47) & convTransposeA_CP_4083_elements(53) & convTransposeA_CP_4083_elements(55);
      gj_convTransposeA_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	83 
    -- CP-element group 57: 	84 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1365/whilex_xbody_ifx_xthen
      -- CP-element group 57: 	 branch_block_stmt_1365/merge_stmt_1746_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1365/merge_stmt_1746__exit__
      -- CP-element group 57: 	 branch_block_stmt_1365/assign_stmt_1752__entry__
      -- CP-element group 57: 	 branch_block_stmt_1365/assign_stmt_1752__exit__
      -- CP-element group 57: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody
      -- CP-element group 57: 	 branch_block_stmt_1365/if_stmt_1740_if_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1365/if_stmt_1740_if_link/if_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1365/assign_stmt_1752/$entry
      -- CP-element group 57: 	 branch_block_stmt_1365/assign_stmt_1752/$exit
      -- CP-element group 57: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/$entry
      -- CP-element group 57: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/$entry
      -- CP-element group 57: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/$entry
      -- CP-element group 57: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/SplitProtocol/$entry
      -- CP-element group 57: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/SplitProtocol/Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/SplitProtocol/Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/SplitProtocol/Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/SplitProtocol/Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1365/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1365/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1365/merge_stmt_1746_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1365/merge_stmt_1746_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1365/merge_stmt_1746_PhiAck/dummy
      -- 
    if_choice_transition_4960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1740_branch_ack_1, ack => convTransposeA_CP_4083_elements(57)); -- 
    rr_5143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(57), ack => type_cast_1639_inst_req_0); -- 
    cr_5148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(57), ack => type_cast_1639_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	62 
    -- CP-element group 58: 	64 
    -- CP-element group 58:  members (24) 
      -- CP-element group 58: 	 branch_block_stmt_1365/whilex_xbody_ifx_xelse
      -- CP-element group 58: 	 branch_block_stmt_1365/merge_stmt_1754__exit__
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796__entry__
      -- CP-element group 58: 	 branch_block_stmt_1365/if_stmt_1740_else_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1365/if_stmt_1740_else_link/else_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/$entry
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1365/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1365/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1365/merge_stmt_1754_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1365/merge_stmt_1754_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1365/merge_stmt_1754_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1365/merge_stmt_1754_PhiAck/dummy
      -- 
    else_choice_transition_4964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1740_branch_ack_0, ack => convTransposeA_CP_4083_elements(58)); -- 
    rr_4980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(58), ack => type_cast_1764_inst_req_0); -- 
    cr_4985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(58), ack => type_cast_1764_inst_req_1); -- 
    cr_4999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(58), ack => type_cast_1773_inst_req_1); -- 
    cr_5013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(58), ack => type_cast_1790_inst_req_1); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_Sample/ra
      -- 
    ra_4981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1764_inst_ack_0, ack => convTransposeA_CP_4083_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1764_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_Sample/rr
      -- 
    ca_4986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1764_inst_ack_1, ack => convTransposeA_CP_4083_elements(60)); -- 
    rr_4994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(60), ack => type_cast_1773_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_Sample/ra
      -- 
    ra_4995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1773_inst_ack_0, ack => convTransposeA_CP_4083_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	58 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1773_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_Sample/rr
      -- 
    ca_5000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1773_inst_ack_1, ack => convTransposeA_CP_4083_elements(62)); -- 
    rr_5008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(62), ack => type_cast_1790_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_Sample/ra
      -- 
    ra_5009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1790_inst_ack_0, ack => convTransposeA_CP_4083_elements(63)); -- 
    -- CP-element group 64:  branch  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	58 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_1365/R_cmp77_1798_place
      -- CP-element group 64: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796__exit__
      -- CP-element group 64: 	 branch_block_stmt_1365/if_stmt_1797__entry__
      -- CP-element group 64: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/$exit
      -- CP-element group 64: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1365/assign_stmt_1760_to_assign_stmt_1796/type_cast_1790_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_1365/if_stmt_1797_dead_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_1365/if_stmt_1797_eval_test/$entry
      -- CP-element group 64: 	 branch_block_stmt_1365/if_stmt_1797_eval_test/$exit
      -- CP-element group 64: 	 branch_block_stmt_1365/if_stmt_1797_eval_test/branch_req
      -- CP-element group 64: 	 branch_block_stmt_1365/if_stmt_1797_if_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_1365/if_stmt_1797_else_link/$entry
      -- 
    ca_5014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1790_inst_ack_1, ack => convTransposeA_CP_4083_elements(64)); -- 
    branch_req_5022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(64), ack => if_stmt_1797_branch_req_0); -- 
    -- CP-element group 65:  merge  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (15) 
      -- CP-element group 65: 	 branch_block_stmt_1365/ifx_xelse_whilex_xend
      -- CP-element group 65: 	 branch_block_stmt_1365/merge_stmt_1803__exit__
      -- CP-element group 65: 	 branch_block_stmt_1365/assign_stmt_1807__entry__
      -- CP-element group 65: 	 branch_block_stmt_1365/if_stmt_1797_if_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1365/if_stmt_1797_if_link/if_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1365/assign_stmt_1807/$entry
      -- CP-element group 65: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1365/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1365/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_1365/merge_stmt_1803_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_1365/merge_stmt_1803_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_1365/merge_stmt_1803_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_1365/merge_stmt_1803_PhiAck/dummy
      -- 
    if_choice_transition_5027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1797_branch_ack_1, ack => convTransposeA_CP_4083_elements(65)); -- 
    req_5044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(65), ack => WPIPE_Block0_done_1805_inst_req_0); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	72 
    -- CP-element group 66: 	73 
    -- CP-element group 66: 	75 
    -- CP-element group 66: 	76 
    -- CP-element group 66:  members (20) 
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 66: 	 branch_block_stmt_1365/if_stmt_1797_else_link/$exit
      -- CP-element group 66: 	 branch_block_stmt_1365/if_stmt_1797_else_link/else_choice_transition
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1797_branch_ack_0, ack => convTransposeA_CP_4083_elements(66)); -- 
    rr_5088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(66), ack => type_cast_1509_inst_req_0); -- 
    cr_5093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(66), ack => type_cast_1509_inst_req_1); -- 
    rr_5111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(66), ack => type_cast_1516_inst_req_0); -- 
    cr_5116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(66), ack => type_cast_1516_inst_req_1); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_update_start_
      -- CP-element group 67: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_Update/req
      -- 
    ack_5045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1805_inst_ack_0, ack => convTransposeA_CP_4083_elements(67)); -- 
    req_5049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(67), ack => WPIPE_Block0_done_1805_inst_req_1); -- 
    -- CP-element group 68:  transition  place  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 branch_block_stmt_1365/$exit
      -- CP-element group 68: 	 branch_block_stmt_1365/branch_block_stmt_1365__exit__
      -- CP-element group 68: 	 branch_block_stmt_1365/assign_stmt_1807__exit__
      -- CP-element group 68: 	 branch_block_stmt_1365/return__
      -- CP-element group 68: 	 branch_block_stmt_1365/merge_stmt_1809__exit__
      -- CP-element group 68: 	 branch_block_stmt_1365/assign_stmt_1807/$exit
      -- CP-element group 68: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1365/assign_stmt_1807/WPIPE_Block0_done_1805_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_1365/return___PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_1365/return___PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_1365/merge_stmt_1809_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_1365/merge_stmt_1809_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_1365/merge_stmt_1809_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_1365/merge_stmt_1809_PhiAck/dummy
      -- 
    ack_5050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1805_inst_ack_1, ack => convTransposeA_CP_4083_elements(68)); -- 
    -- CP-element group 69:  transition  output  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	29 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/$exit
      -- CP-element group 69: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1507_konst_delay_trans
      -- CP-element group 69: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_req
      -- 
    phi_stmt_1503_req_5061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1503_req_5061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(69), ack => phi_stmt_1503_req_0); -- 
    -- Element group convTransposeA_CP_4083_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => convTransposeA_CP_4083_elements(29), ack => convTransposeA_CP_4083_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  transition  output  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/$exit
      -- CP-element group 70: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1514_konst_delay_trans
      -- CP-element group 70: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_req
      -- 
    phi_stmt_1510_req_5069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1510_req_5069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(70), ack => phi_stmt_1510_req_0); -- 
    -- Element group convTransposeA_CP_4083_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convTransposeA_CP_4083_elements(29), ack => convTransposeA_CP_4083_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	79 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1365/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(69) & convTransposeA_CP_4083_elements(70);
      gj_convTransposeA_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	66 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/SplitProtocol/Sample/ra
      -- 
    ra_5089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1509_inst_ack_0, ack => convTransposeA_CP_4083_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	66 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/SplitProtocol/Update/ca
      -- 
    ca_5094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1509_inst_ack_1, ack => convTransposeA_CP_4083_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	78 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/$exit
      -- CP-element group 74: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/$exit
      -- CP-element group 74: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_sources/type_cast_1509/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1503/phi_stmt_1503_req
      -- 
    phi_stmt_1503_req_5095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1503_req_5095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(74), ack => phi_stmt_1503_req_1); -- 
    convTransposeA_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(72) & convTransposeA_CP_4083_elements(73);
      gj_convTransposeA_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	66 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/SplitProtocol/Sample/ra
      -- 
    ra_5112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1516_inst_ack_0, ack => convTransposeA_CP_4083_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	66 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/SplitProtocol/Update/ca
      -- 
    ca_5117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1516_inst_ack_1, ack => convTransposeA_CP_4083_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/$exit
      -- CP-element group 77: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/$exit
      -- CP-element group 77: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_sources/type_cast_1516/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1510/phi_stmt_1510_req
      -- 
    phi_stmt_1510_req_5118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1510_req_5118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(77), ack => phi_stmt_1510_req_1); -- 
    convTransposeA_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(75) & convTransposeA_CP_4083_elements(76);
      gj_convTransposeA_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	74 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1365/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(74) & convTransposeA_CP_4083_elements(77);
      gj_convTransposeA_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  merge  fork  transition  place  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	71 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1365/merge_stmt_1502_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_1365/merge_stmt_1502_PhiAck/$entry
      -- 
    convTransposeA_CP_4083_elements(79) <= OrReduce(convTransposeA_CP_4083_elements(71) & convTransposeA_CP_4083_elements(78));
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1365/merge_stmt_1502_PhiAck/phi_stmt_1503_ack
      -- 
    phi_stmt_1503_ack_5123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1503_ack_0, ack => convTransposeA_CP_4083_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1365/merge_stmt_1502_PhiAck/phi_stmt_1510_ack
      -- 
    phi_stmt_1510_ack_5124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1510_ack_0, ack => convTransposeA_CP_4083_elements(81)); -- 
    -- CP-element group 82:  join  fork  transition  place  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	31 
    -- CP-element group 82: 	32 
    -- CP-element group 82: 	33 
    -- CP-element group 82: 	30 
    -- CP-element group 82:  members (16) 
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1365/merge_stmt_1502__exit__
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630__entry__
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/$entry
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1527_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_1365/assign_stmt_1523_to_assign_stmt_1630/type_cast_1522_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1365/merge_stmt_1502_PhiAck/$exit
      -- 
    cr_4695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(82), ack => type_cast_1527_inst_req_1); -- 
    rr_4690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(82), ack => type_cast_1527_inst_req_0); -- 
    cr_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(82), ack => type_cast_1522_inst_req_1); -- 
    rr_4676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(82), ack => type_cast_1522_inst_req_0); -- 
    convTransposeA_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(80) & convTransposeA_CP_4083_elements(81);
      gj_convTransposeA_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	57 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/SplitProtocol/Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/SplitProtocol/Sample/ra
      -- 
    ra_5144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1639_inst_ack_0, ack => convTransposeA_CP_4083_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	57 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/SplitProtocol/Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/SplitProtocol/Update/ca
      -- 
    ca_5149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1639_inst_ack_1, ack => convTransposeA_CP_4083_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/$exit
      -- CP-element group 85: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/$exit
      -- CP-element group 85: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1639/SplitProtocol/$exit
      -- CP-element group 85: 	 branch_block_stmt_1365/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_req
      -- 
    phi_stmt_1633_req_5150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1633_req_5150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(85), ack => phi_stmt_1633_req_1); -- 
    convTransposeA_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(83) & convTransposeA_CP_4083_elements(84);
      gj_convTransposeA_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  output  delay-element  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	34 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1365/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_1365/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1633/$exit
      -- CP-element group 86: 	 branch_block_stmt_1365/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1365/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_sources/type_cast_1637_konst_delay_trans
      -- CP-element group 86: 	 branch_block_stmt_1365/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1633/phi_stmt_1633_req
      -- 
    phi_stmt_1633_req_5161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1633_req_5161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(86), ack => phi_stmt_1633_req_0); -- 
    -- Element group convTransposeA_CP_4083_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => convTransposeA_CP_4083_elements(34), ack => convTransposeA_CP_4083_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  merge  transition  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1365/merge_stmt_1632_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_1365/merge_stmt_1632_PhiAck/$entry
      -- 
    convTransposeA_CP_4083_elements(87) <= OrReduce(convTransposeA_CP_4083_elements(85) & convTransposeA_CP_4083_elements(86));
    -- CP-element group 88:  fork  transition  place  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	35 
    -- CP-element group 88: 	36 
    -- CP-element group 88: 	38 
    -- CP-element group 88: 	40 
    -- CP-element group 88: 	42 
    -- CP-element group 88: 	44 
    -- CP-element group 88: 	46 
    -- CP-element group 88: 	48 
    -- CP-element group 88: 	50 
    -- CP-element group 88: 	53 
    -- CP-element group 88: 	54 
    -- CP-element group 88: 	55 
    -- CP-element group 88:  members (45) 
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1687_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1711_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/merge_stmt_1632__exit__
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739__entry__
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1680_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1691_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1649_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1686_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/array_obj_ref_1717_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/addr_of_1718_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/ptr_deref_1721_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1365/assign_stmt_1646_to_assign_stmt_1739/type_cast_1727_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1365/merge_stmt_1632_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_1365/merge_stmt_1632_PhiAck/phi_stmt_1633_ack
      -- 
    phi_stmt_1633_ack_5166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1633_ack_0, ack => convTransposeA_CP_4083_elements(88)); -- 
    req_4772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => addr_of_1687_final_reg_req_1); -- 
    cr_4817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => ptr_deref_1691_load_0_req_1); -- 
    cr_4726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1680_inst_req_1); -- 
    cr_4836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1711_inst_req_1); -- 
    req_4757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => array_obj_ref_1686_index_offset_req_1); -- 
    cr_4712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1649_inst_req_1); -- 
    rr_4707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1649_inst_req_0); -- 
    req_4867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => array_obj_ref_1717_index_offset_req_1); -- 
    req_4882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => addr_of_1718_final_reg_req_1); -- 
    cr_4932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => ptr_deref_1721_store_0_req_1); -- 
    rr_4941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1727_inst_req_0); -- 
    cr_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1727_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1592_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1613_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1673_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1705_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1421_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1421_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom52_1716_resized : std_logic_vector(13 downto 0);
    signal R_idxprom52_1716_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1685_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1685_scaled : std_logic_vector(13 downto 0);
    signal add16_1553 : std_logic_vector(31 downto 0);
    signal add27_1568 : std_logic_vector(31 downto 0);
    signal add42_1625 : std_logic_vector(31 downto 0);
    signal add44_1660 : std_logic_vector(31 downto 0);
    signal add57_1734 : std_logic_vector(31 downto 0);
    signal add8_1655 : std_logic_vector(31 downto 0);
    signal add_1538 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1686_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1686_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1717_root_address : std_logic_vector(13 downto 0);
    signal arrayidx53_1719 : std_logic_vector(31 downto 0);
    signal arrayidx_1688 : std_logic_vector(31 downto 0);
    signal call_1368 : std_logic_vector(15 downto 0);
    signal cmp68_1770 : std_logic_vector(0 downto 0);
    signal cmp77_1796 : std_logic_vector(0 downto 0);
    signal cmp_1739 : std_logic_vector(0 downto 0);
    signal conv13_1407 : std_logic_vector(31 downto 0);
    signal conv18_1426 : std_logic_vector(31 downto 0);
    signal conv24_1440 : std_logic_vector(31 downto 0);
    signal conv37_1594 : std_logic_vector(31 downto 0);
    signal conv3_1523 : std_logic_vector(31 downto 0);
    signal conv40_1615 : std_logic_vector(31 downto 0);
    signal conv56_1728 : std_logic_vector(31 downto 0);
    signal conv66_1765 : std_logic_vector(31 downto 0);
    signal conv6_1528 : std_logic_vector(31 downto 0);
    signal conv74_1791 : std_logic_vector(31 downto 0);
    signal conv90_1650 : std_logic_vector(31 downto 0);
    signal div76_1500 : std_logic_vector(31 downto 0);
    signal div_1482 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1490 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1377 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1389 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1399 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1415 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1432 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1448 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1460 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1472 : std_logic_vector(31 downto 0);
    signal idxprom52_1712 : std_logic_vector(63 downto 0);
    signal idxprom_1681 : std_logic_vector(63 downto 0);
    signal inc72_1774 : std_logic_vector(15 downto 0);
    signal inc72x_xinput_dim0x_x2_1779 : std_logic_vector(15 downto 0);
    signal inc_1760 : std_logic_vector(15 downto 0);
    signal indvar_1633 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1752 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1510 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1503 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1786 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1646 : std_logic_vector(15 downto 0);
    signal mul14_1548 : std_logic_vector(31 downto 0);
    signal mul25_1563 : std_logic_vector(31 downto 0);
    signal mul41_1620 : std_logic_vector(31 downto 0);
    signal mul43_1630 : std_logic_vector(31 downto 0);
    signal mul7_1543 : std_logic_vector(31 downto 0);
    signal mul_1533 : std_logic_vector(31 downto 0);
    signal ptr_deref_1380_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1380_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1380_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1380_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1380_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1392_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1392_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1392_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1392_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1392_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1402_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1402_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1402_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1402_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1402_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1418_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1418_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1418_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1418_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1418_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1435_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1435_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1435_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1435_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1435_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1451_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1451_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1451_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1451_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1451_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1463_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1463_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1463_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1463_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1463_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1475_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1475_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1475_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1475_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1475_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1493_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1493_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1493_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1493_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1493_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1691_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1691_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1691_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1691_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1691_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1721_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1721_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1721_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1721_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1721_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1721_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext91_1606 : std_logic_vector(31 downto 0);
    signal sext93_1666 : std_logic_vector(31 downto 0);
    signal sext94_1698 : std_logic_vector(31 downto 0);
    signal sext_1585 : std_logic_vector(31 downto 0);
    signal shr51_1707 : std_logic_vector(31 downto 0);
    signal shr_1675 : std_logic_vector(31 downto 0);
    signal sub19_1600 : std_logic_vector(31 downto 0);
    signal sub30_1573 : std_logic_vector(31 downto 0);
    signal sub31_1579 : std_logic_vector(31 downto 0);
    signal sub_1558 : std_logic_vector(31 downto 0);
    signal tmp12_1403 : std_logic_vector(15 downto 0);
    signal tmp15_1419 : std_logic_vector(31 downto 0);
    signal tmp17_1422 : std_logic_vector(15 downto 0);
    signal tmp1_1381 : std_logic_vector(31 downto 0);
    signal tmp23_1436 : std_logic_vector(15 downto 0);
    signal tmp26_1452 : std_logic_vector(31 downto 0);
    signal tmp35_1464 : std_logic_vector(31 downto 0);
    signal tmp38_1476 : std_logic_vector(31 downto 0);
    signal tmp48_1692 : std_logic_vector(63 downto 0);
    signal tmp4_1393 : std_logic_vector(31 downto 0);
    signal tmp75_1494 : std_logic_vector(31 downto 0);
    signal type_cast_1480_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1498_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1507_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1509_wire : std_logic_vector(15 downto 0);
    signal type_cast_1514_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1516_wire : std_logic_vector(15 downto 0);
    signal type_cast_1521_wire : std_logic_vector(31 downto 0);
    signal type_cast_1526_wire : std_logic_vector(31 downto 0);
    signal type_cast_1577_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1583_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1588_wire : std_logic_vector(31 downto 0);
    signal type_cast_1591_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1598_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1604_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1609_wire : std_logic_vector(31 downto 0);
    signal type_cast_1612_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1637_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1639_wire : std_logic_vector(15 downto 0);
    signal type_cast_1644_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1664_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1669_wire : std_logic_vector(31 downto 0);
    signal type_cast_1672_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1679_wire : std_logic_vector(63 downto 0);
    signal type_cast_1696_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1701_wire : std_logic_vector(31 downto 0);
    signal type_cast_1704_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1710_wire : std_logic_vector(63 downto 0);
    signal type_cast_1726_wire : std_logic_vector(31 downto 0);
    signal type_cast_1732_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1750_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1758_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1763_wire : std_logic_vector(31 downto 0);
    signal type_cast_1783_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1789_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1421_word_address_0 <= "0";
    array_obj_ref_1686_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1686_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1686_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1686_resized_base_address <= "00000000000000";
    array_obj_ref_1717_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1717_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1717_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1717_resized_base_address <= "00000000000000";
    iNsTr_10_1490 <= "00000000000000000000000000000010";
    iNsTr_2_1377 <= "00000000000000000000000000000100";
    iNsTr_3_1389 <= "00000000000000000000000000000011";
    iNsTr_4_1399 <= "00000000000000000000000000000000";
    iNsTr_5_1415 <= "00000000000000000000000000000011";
    iNsTr_6_1432 <= "00000000000000000000000000000001";
    iNsTr_7_1448 <= "00000000000000000000000000000100";
    iNsTr_8_1460 <= "00000000000000000000000000000100";
    iNsTr_9_1472 <= "00000000000000000000000000000011";
    ptr_deref_1380_word_offset_0 <= "0000000";
    ptr_deref_1392_word_offset_0 <= "0000000";
    ptr_deref_1402_word_offset_0 <= "0";
    ptr_deref_1418_word_offset_0 <= "0000000";
    ptr_deref_1435_word_offset_0 <= "0";
    ptr_deref_1451_word_offset_0 <= "0000000";
    ptr_deref_1463_word_offset_0 <= "0000000";
    ptr_deref_1475_word_offset_0 <= "0000000";
    ptr_deref_1493_word_offset_0 <= "0000000";
    ptr_deref_1691_word_offset_0 <= "00000000000000";
    ptr_deref_1721_word_offset_0 <= "00000000000000";
    type_cast_1480_wire_constant <= "00000000000000000000000000000001";
    type_cast_1498_wire_constant <= "00000000000000000000000000000001";
    type_cast_1507_wire_constant <= "0000000000000000";
    type_cast_1514_wire_constant <= "0000000000000000";
    type_cast_1577_wire_constant <= "00000000000000000000000000010000";
    type_cast_1583_wire_constant <= "11111111111111110000000000000000";
    type_cast_1591_wire_constant <= "00000000000000000000000000010000";
    type_cast_1598_wire_constant <= "00000000000000000000000000010000";
    type_cast_1604_wire_constant <= "11111111111111110000000000000000";
    type_cast_1612_wire_constant <= "00000000000000000000000000010000";
    type_cast_1637_wire_constant <= "0000000000000000";
    type_cast_1644_wire_constant <= "0000000000000100";
    type_cast_1664_wire_constant <= "00000000000000000000000000010000";
    type_cast_1672_wire_constant <= "00000000000000000000000000010010";
    type_cast_1696_wire_constant <= "00000000000000000000000000010000";
    type_cast_1704_wire_constant <= "00000000000000000000000000010010";
    type_cast_1732_wire_constant <= "00000000000000000000000000000100";
    type_cast_1750_wire_constant <= "0000000000000001";
    type_cast_1758_wire_constant <= "0000000000000001";
    type_cast_1783_wire_constant <= "0000000000000000";
    phi_stmt_1503: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1507_wire_constant & type_cast_1509_wire;
      req <= phi_stmt_1503_req_0 & phi_stmt_1503_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1503",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1503_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1503,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1503
    phi_stmt_1510: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1514_wire_constant & type_cast_1516_wire;
      req <= phi_stmt_1510_req_0 & phi_stmt_1510_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1510",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1510_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1510,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1510
    phi_stmt_1633: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1637_wire_constant & type_cast_1639_wire;
      req <= phi_stmt_1633_req_0 & phi_stmt_1633_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1633",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1633_ack_0,
          idata => idata,
          odata => indvar_1633,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1633
    -- flow-through select operator MUX_1785_inst
    input_dim1x_x2_1786 <= type_cast_1783_wire_constant when (cmp68_1770(0) /=  '0') else inc_1760;
    addr_of_1687_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1687_final_reg_req_0;
      addr_of_1687_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1687_final_reg_req_1;
      addr_of_1687_final_reg_ack_1<= rack(0);
      addr_of_1687_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1687_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1686_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1688,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1718_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1718_final_reg_req_0;
      addr_of_1718_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1718_final_reg_req_1;
      addr_of_1718_final_reg_ack_1<= rack(0);
      addr_of_1718_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1718_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1717_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx53_1719,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1406_inst_req_0;
      type_cast_1406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1406_inst_req_1;
      type_cast_1406_inst_ack_1<= rack(0);
      type_cast_1406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_1403,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_1407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1425_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1425_inst_req_0;
      type_cast_1425_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1425_inst_req_1;
      type_cast_1425_inst_ack_1<= rack(0);
      type_cast_1425_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1425_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp17_1422,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_1426,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1439_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1439_inst_req_0;
      type_cast_1439_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1439_inst_req_1;
      type_cast_1439_inst_ack_1<= rack(0);
      type_cast_1439_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1439_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp23_1436,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_1440,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1509_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1509_inst_req_0;
      type_cast_1509_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1509_inst_req_1;
      type_cast_1509_inst_ack_1<= rack(0);
      type_cast_1509_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1509_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1509_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1516_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1516_inst_req_0;
      type_cast_1516_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1516_inst_req_1;
      type_cast_1516_inst_ack_1<= rack(0);
      type_cast_1516_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1516_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc72x_xinput_dim0x_x2_1779,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1516_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1522_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1522_inst_req_0;
      type_cast_1522_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1522_inst_req_1;
      type_cast_1522_inst_ack_1<= rack(0);
      type_cast_1522_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1522_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1521_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1523,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1527_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1527_inst_req_0;
      type_cast_1527_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1527_inst_req_1;
      type_cast_1527_inst_ack_1<= rack(0);
      type_cast_1527_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1527_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1526_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv6_1528,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1588_inst
    process(sext_1585) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_1585(31 downto 0);
      type_cast_1588_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1593_inst
    process(ASHR_i32_i32_1592_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1592_wire(31 downto 0);
      conv37_1594 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1609_inst
    process(sext91_1606) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext91_1606(31 downto 0);
      type_cast_1609_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1614_inst
    process(ASHR_i32_i32_1613_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1613_wire(31 downto 0);
      conv40_1615 <= tmp_var; -- 
    end process;
    type_cast_1639_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1639_inst_req_0;
      type_cast_1639_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1639_inst_req_1;
      type_cast_1639_inst_ack_1<= rack(0);
      type_cast_1639_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1639_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1752,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1639_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1649_inst_req_0;
      type_cast_1649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1649_inst_req_1;
      type_cast_1649_inst_ack_1<= rack(0);
      type_cast_1649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1669_inst
    process(sext93_1666) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext93_1666(31 downto 0);
      type_cast_1669_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1674_inst
    process(ASHR_i32_i32_1673_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1673_wire(31 downto 0);
      shr_1675 <= tmp_var; -- 
    end process;
    type_cast_1680_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1680_inst_req_0;
      type_cast_1680_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1680_inst_req_1;
      type_cast_1680_inst_ack_1<= rack(0);
      type_cast_1680_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1680_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1679_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1681,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1701_inst
    process(sext94_1698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext94_1698(31 downto 0);
      type_cast_1701_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1706_inst
    process(ASHR_i32_i32_1705_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1705_wire(31 downto 0);
      shr51_1707 <= tmp_var; -- 
    end process;
    type_cast_1711_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1711_inst_req_0;
      type_cast_1711_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1711_inst_req_1;
      type_cast_1711_inst_ack_1<= rack(0);
      type_cast_1711_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1711_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1710_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom52_1712,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1727_inst_req_0;
      type_cast_1727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1727_inst_req_1;
      type_cast_1727_inst_ack_1<= rack(0);
      type_cast_1727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1726_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_1728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1764_inst_req_0;
      type_cast_1764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1764_inst_req_1;
      type_cast_1764_inst_ack_1<= rack(0);
      type_cast_1764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1763_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1773_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1773_inst_req_0;
      type_cast_1773_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1773_inst_req_1;
      type_cast_1773_inst_ack_1<= rack(0);
      type_cast_1773_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1773_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp68_1770,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc72_1774,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1790_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1790_inst_req_0;
      type_cast_1790_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1790_inst_req_1;
      type_cast_1790_inst_ack_1<= rack(0);
      type_cast_1790_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1790_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1789_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_1791,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1421_gather_scatter
    process(LOAD_padding_1421_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1421_data_0;
      ov(15 downto 0) := iv;
      tmp17_1422 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1686_index_1_rename
    process(R_idxprom_1685_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1685_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1685_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1686_index_1_resize
    process(idxprom_1681) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1681;
      ov := iv(13 downto 0);
      R_idxprom_1685_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1686_root_address_inst
    process(array_obj_ref_1686_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1686_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1686_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1717_index_1_rename
    process(R_idxprom52_1716_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom52_1716_resized;
      ov(13 downto 0) := iv;
      R_idxprom52_1716_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1717_index_1_resize
    process(idxprom52_1712) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom52_1712;
      ov := iv(13 downto 0);
      R_idxprom52_1716_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1717_root_address_inst
    process(array_obj_ref_1717_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1717_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1717_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1380_addr_0
    process(ptr_deref_1380_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1380_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1380_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1380_base_resize
    process(iNsTr_2_1377) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1377;
      ov := iv(6 downto 0);
      ptr_deref_1380_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1380_gather_scatter
    process(ptr_deref_1380_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1380_data_0;
      ov(31 downto 0) := iv;
      tmp1_1381 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1380_root_address_inst
    process(ptr_deref_1380_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1380_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1380_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1392_addr_0
    process(ptr_deref_1392_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1392_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1392_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1392_base_resize
    process(iNsTr_3_1389) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1389;
      ov := iv(6 downto 0);
      ptr_deref_1392_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1392_gather_scatter
    process(ptr_deref_1392_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1392_data_0;
      ov(31 downto 0) := iv;
      tmp4_1393 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1392_root_address_inst
    process(ptr_deref_1392_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1392_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1392_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1402_addr_0
    process(ptr_deref_1402_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1402_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1402_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1402_base_resize
    process(iNsTr_4_1399) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1399;
      ov := iv(0 downto 0);
      ptr_deref_1402_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1402_gather_scatter
    process(ptr_deref_1402_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1402_data_0;
      ov(15 downto 0) := iv;
      tmp12_1403 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1402_root_address_inst
    process(ptr_deref_1402_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1402_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1402_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1418_addr_0
    process(ptr_deref_1418_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1418_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1418_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1418_base_resize
    process(iNsTr_5_1415) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1415;
      ov := iv(6 downto 0);
      ptr_deref_1418_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1418_gather_scatter
    process(ptr_deref_1418_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1418_data_0;
      ov(31 downto 0) := iv;
      tmp15_1419 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1418_root_address_inst
    process(ptr_deref_1418_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1418_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1418_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1435_addr_0
    process(ptr_deref_1435_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1435_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1435_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1435_base_resize
    process(iNsTr_6_1432) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1432;
      ov := iv(0 downto 0);
      ptr_deref_1435_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1435_gather_scatter
    process(ptr_deref_1435_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1435_data_0;
      ov(15 downto 0) := iv;
      tmp23_1436 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1435_root_address_inst
    process(ptr_deref_1435_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1435_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1435_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1451_addr_0
    process(ptr_deref_1451_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1451_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1451_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1451_base_resize
    process(iNsTr_7_1448) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1448;
      ov := iv(6 downto 0);
      ptr_deref_1451_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1451_gather_scatter
    process(ptr_deref_1451_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1451_data_0;
      ov(31 downto 0) := iv;
      tmp26_1452 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1451_root_address_inst
    process(ptr_deref_1451_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1451_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1451_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1463_addr_0
    process(ptr_deref_1463_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1463_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1463_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1463_base_resize
    process(iNsTr_8_1460) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1460;
      ov := iv(6 downto 0);
      ptr_deref_1463_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1463_gather_scatter
    process(ptr_deref_1463_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1463_data_0;
      ov(31 downto 0) := iv;
      tmp35_1464 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1463_root_address_inst
    process(ptr_deref_1463_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1463_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1463_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1475_addr_0
    process(ptr_deref_1475_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1475_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1475_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1475_base_resize
    process(iNsTr_9_1472) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1472;
      ov := iv(6 downto 0);
      ptr_deref_1475_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1475_gather_scatter
    process(ptr_deref_1475_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1475_data_0;
      ov(31 downto 0) := iv;
      tmp38_1476 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1475_root_address_inst
    process(ptr_deref_1475_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1475_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1475_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1493_addr_0
    process(ptr_deref_1493_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1493_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1493_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1493_base_resize
    process(iNsTr_10_1490) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1490;
      ov := iv(6 downto 0);
      ptr_deref_1493_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1493_gather_scatter
    process(ptr_deref_1493_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1493_data_0;
      ov(31 downto 0) := iv;
      tmp75_1494 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1493_root_address_inst
    process(ptr_deref_1493_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1493_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1493_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1691_addr_0
    process(ptr_deref_1691_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1691_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1691_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1691_base_resize
    process(arrayidx_1688) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1688;
      ov := iv(13 downto 0);
      ptr_deref_1691_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1691_gather_scatter
    process(ptr_deref_1691_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1691_data_0;
      ov(63 downto 0) := iv;
      tmp48_1692 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1691_root_address_inst
    process(ptr_deref_1691_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1691_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1691_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1721_addr_0
    process(ptr_deref_1721_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1721_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1721_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1721_base_resize
    process(arrayidx53_1719) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx53_1719;
      ov := iv(13 downto 0);
      ptr_deref_1721_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1721_gather_scatter
    process(tmp48_1692) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp48_1692;
      ov(63 downto 0) := iv;
      ptr_deref_1721_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1721_root_address_inst
    process(ptr_deref_1721_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1721_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1721_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1740_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1739;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1740_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1740_branch_req_0,
          ack0 => if_stmt_1740_branch_ack_0,
          ack1 => if_stmt_1740_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1797_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_1796;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1797_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1797_branch_req_0,
          ack0 => if_stmt_1797_branch_ack_0,
          ack1 => if_stmt_1797_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1751_inst
    process(indvar_1633) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1633, type_cast_1750_wire_constant, tmp_var);
      indvarx_xnext_1752 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1759_inst
    process(input_dim1x_x1x_xph_1503) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1503, type_cast_1758_wire_constant, tmp_var);
      inc_1760 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1778_inst
    process(inc72_1774, input_dim0x_x2x_xph_1510) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc72_1774, input_dim0x_x2x_xph_1510, tmp_var);
      inc72x_xinput_dim0x_x2_1779 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1537_inst
    process(mul_1533, conv3_1523) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_1533, conv3_1523, tmp_var);
      add_1538 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1552_inst
    process(mul14_1548, tmp15_1419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul14_1548, tmp15_1419, tmp_var);
      add16_1553 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1567_inst
    process(mul25_1563, tmp26_1452) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul25_1563, tmp26_1452, tmp_var);
      add27_1568 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1584_inst
    process(sub31_1579) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub31_1579, type_cast_1583_wire_constant, tmp_var);
      sext_1585 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1605_inst
    process(sub19_1600) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub19_1600, type_cast_1604_wire_constant, tmp_var);
      sext91_1606 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1624_inst
    process(conv37_1594, mul41_1620) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv37_1594, mul41_1620, tmp_var);
      add42_1625 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1654_inst
    process(mul7_1543, conv90_1650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul7_1543, conv90_1650, tmp_var);
      add8_1655 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1659_inst
    process(mul43_1630, conv90_1650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul43_1630, conv90_1650, tmp_var);
      add44_1660 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1733_inst
    process(conv56_1728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv56_1728, type_cast_1732_wire_constant, tmp_var);
      add57_1734 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1592_inst
    process(type_cast_1588_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1588_wire, type_cast_1591_wire_constant, tmp_var);
      ASHR_i32_i32_1592_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1613_inst
    process(type_cast_1609_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1609_wire, type_cast_1612_wire_constant, tmp_var);
      ASHR_i32_i32_1613_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1673_inst
    process(type_cast_1669_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1669_wire, type_cast_1672_wire_constant, tmp_var);
      ASHR_i32_i32_1673_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1705_inst
    process(type_cast_1701_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1701_wire, type_cast_1704_wire_constant, tmp_var);
      ASHR_i32_i32_1705_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1769_inst
    process(conv66_1765, div_1482) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv66_1765, div_1482, tmp_var);
      cmp68_1770 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1795_inst
    process(conv74_1791, div76_1500) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv74_1791, div76_1500, tmp_var);
      cmp77_1796 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1481_inst
    process(tmp4_1393) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1393, type_cast_1480_wire_constant, tmp_var);
      div_1482 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1499_inst
    process(tmp75_1494) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp75_1494, type_cast_1498_wire_constant, tmp_var);
      div76_1500 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1645_inst
    process(indvar_1633) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1633, type_cast_1644_wire_constant, tmp_var);
      input_dim2x_x1_1646 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1532_inst
    process(tmp4_1393, conv6_1528) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp4_1393, conv6_1528, tmp_var);
      mul_1533 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1542_inst
    process(add_1538, tmp1_1381) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1538, tmp1_1381, tmp_var);
      mul7_1543 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1547_inst
    process(conv13_1407, conv6_1528) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv13_1407, conv6_1528, tmp_var);
      mul14_1548 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1562_inst
    process(conv24_1440, conv3_1523) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv24_1440, conv3_1523, tmp_var);
      mul25_1563 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1619_inst
    process(tmp38_1476, conv40_1615) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp38_1476, conv40_1615, tmp_var);
      mul41_1620 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1629_inst
    process(add42_1625, tmp35_1464) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add42_1625, tmp35_1464, tmp_var);
      mul43_1630 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1578_inst
    process(sub30_1573) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub30_1573, type_cast_1577_wire_constant, tmp_var);
      sub31_1579 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1599_inst
    process(sub_1558) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_1558, type_cast_1598_wire_constant, tmp_var);
      sub19_1600 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1665_inst
    process(add8_1655) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add8_1655, type_cast_1664_wire_constant, tmp_var);
      sext93_1666 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1697_inst
    process(add44_1660) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add44_1660, type_cast_1696_wire_constant, tmp_var);
      sext94_1698 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1557_inst
    process(add16_1553, conv18_1426) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add16_1553, conv18_1426, tmp_var);
      sub_1558 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1572_inst
    process(add27_1568, conv18_1426) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add27_1568, conv18_1426, tmp_var);
      sub30_1573 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1738_inst
    process(add57_1734, tmp1_1381) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add57_1734, tmp1_1381, tmp_var);
      cmp_1739 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_1686_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1685_scaled;
      array_obj_ref_1686_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1686_index_offset_req_0;
      array_obj_ref_1686_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1686_index_offset_req_1;
      array_obj_ref_1686_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_1717_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom52_1716_scaled;
      array_obj_ref_1717_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1717_index_offset_req_0;
      array_obj_ref_1717_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1717_index_offset_req_1;
      array_obj_ref_1717_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- unary operator type_cast_1521_inst
    process(input_dim1x_x1x_xph_1503) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_1503, tmp_var);
      type_cast_1521_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1526_inst
    process(input_dim0x_x2x_xph_1510) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_1510, tmp_var);
      type_cast_1526_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1679_inst
    process(shr_1675) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1675, tmp_var);
      type_cast_1679_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1710_inst
    process(shr51_1707) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr51_1707, tmp_var);
      type_cast_1710_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1726_inst
    process(input_dim2x_x1_1646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1646, tmp_var);
      type_cast_1726_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1763_inst
    process(inc_1760) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1760, tmp_var);
      type_cast_1763_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1789_inst
    process(inc72x_xinput_dim0x_x2_1779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc72x_xinput_dim0x_x2_1779, tmp_var);
      type_cast_1789_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1421_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1421_load_0_req_0;
      LOAD_padding_1421_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1421_load_0_req_1;
      LOAD_padding_1421_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1421_word_address_0;
      LOAD_padding_1421_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1493_load_0 ptr_deref_1380_load_0 ptr_deref_1392_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1493_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1380_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1392_load_0_req_0;
      ptr_deref_1493_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1380_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1392_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1493_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1380_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1392_load_0_req_1;
      ptr_deref_1493_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1380_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1392_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1493_word_address_0 & ptr_deref_1380_word_address_0 & ptr_deref_1392_word_address_0;
      ptr_deref_1493_data_0 <= data_out(95 downto 64);
      ptr_deref_1380_data_0 <= data_out(63 downto 32);
      ptr_deref_1392_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1435_load_0 ptr_deref_1402_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1435_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1402_load_0_req_0;
      ptr_deref_1435_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1402_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1435_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1402_load_0_req_1;
      ptr_deref_1435_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1402_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1435_word_address_0 & ptr_deref_1402_word_address_0;
      ptr_deref_1435_data_0 <= data_out(31 downto 16);
      ptr_deref_1402_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1451_load_0 ptr_deref_1418_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1451_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1418_load_0_req_0;
      ptr_deref_1451_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1418_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1451_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1418_load_0_req_1;
      ptr_deref_1451_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1418_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1451_word_address_0 & ptr_deref_1418_word_address_0;
      ptr_deref_1451_data_0 <= data_out(63 downto 32);
      ptr_deref_1418_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1463_load_0 ptr_deref_1475_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1463_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1475_load_0_req_0;
      ptr_deref_1463_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1475_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1463_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1475_load_0_req_1;
      ptr_deref_1463_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1475_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1463_word_address_0 & ptr_deref_1475_word_address_0;
      ptr_deref_1463_data_0 <= data_out(63 downto 32);
      ptr_deref_1475_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1691_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1691_load_0_req_0;
      ptr_deref_1691_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1691_load_0_req_1;
      ptr_deref_1691_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1691_word_address_0;
      ptr_deref_1691_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_1721_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1721_store_0_req_0;
      ptr_deref_1721_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1721_store_0_req_1;
      ptr_deref_1721_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1721_word_address_0;
      data_in <= ptr_deref_1721_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1367_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_start_1367_inst_req_0;
      RPIPE_Block0_start_1367_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_start_1367_inst_req_1;
      RPIPE_Block0_start_1367_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1368 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1805_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1805_inst_req_0;
      WPIPE_Block0_done_1805_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1805_inst_req_1;
      WPIPE_Block0_done_1805_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1368;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_5207_start: Boolean;
  signal convTransposeB_CP_5207_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1864_inst_ack_0 : boolean;
  signal type_cast_1864_inst_req_0 : boolean;
  signal type_cast_1883_inst_req_1 : boolean;
  signal type_cast_1883_inst_ack_1 : boolean;
  signal ptr_deref_1909_load_0_req_0 : boolean;
  signal ptr_deref_1909_load_0_ack_1 : boolean;
  signal ptr_deref_1909_load_0_ack_0 : boolean;
  signal LOAD_padding_1879_load_0_req_1 : boolean;
  signal ptr_deref_1909_load_0_req_1 : boolean;
  signal type_cast_1897_inst_req_0 : boolean;
  signal type_cast_1897_inst_ack_0 : boolean;
  signal LOAD_padding_1879_load_0_ack_1 : boolean;
  signal ptr_deref_1876_load_0_ack_1 : boolean;
  signal type_cast_1897_inst_req_1 : boolean;
  signal type_cast_1897_inst_ack_1 : boolean;
  signal ptr_deref_1893_load_0_req_1 : boolean;
  signal ptr_deref_1893_load_0_ack_1 : boolean;
  signal type_cast_1883_inst_req_0 : boolean;
  signal type_cast_1883_inst_ack_0 : boolean;
  signal type_cast_1864_inst_req_1 : boolean;
  signal ptr_deref_1876_load_0_req_1 : boolean;
  signal LOAD_padding_1879_load_0_req_0 : boolean;
  signal LOAD_padding_1879_load_0_ack_0 : boolean;
  signal ptr_deref_1876_load_0_req_0 : boolean;
  signal ptr_deref_1921_load_0_req_1 : boolean;
  signal ptr_deref_1921_load_0_ack_1 : boolean;
  signal ptr_deref_1893_load_0_req_0 : boolean;
  signal ptr_deref_1893_load_0_ack_0 : boolean;
  signal ptr_deref_1876_load_0_ack_0 : boolean;
  signal ptr_deref_1921_load_0_req_0 : boolean;
  signal ptr_deref_1921_load_0_ack_0 : boolean;
  signal type_cast_1864_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1815_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1815_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1815_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1815_inst_ack_1 : boolean;
  signal ptr_deref_1828_load_0_req_0 : boolean;
  signal ptr_deref_1828_load_0_ack_0 : boolean;
  signal ptr_deref_1828_load_0_req_1 : boolean;
  signal ptr_deref_1828_load_0_ack_1 : boolean;
  signal type_cast_1838_inst_req_0 : boolean;
  signal type_cast_1838_inst_ack_0 : boolean;
  signal type_cast_1838_inst_req_1 : boolean;
  signal type_cast_1838_inst_ack_1 : boolean;
  signal ptr_deref_1850_load_0_req_0 : boolean;
  signal ptr_deref_1850_load_0_ack_0 : boolean;
  signal ptr_deref_1850_load_0_req_1 : boolean;
  signal ptr_deref_1850_load_0_ack_1 : boolean;
  signal ptr_deref_1860_load_0_req_0 : boolean;
  signal ptr_deref_1860_load_0_ack_0 : boolean;
  signal ptr_deref_1860_load_0_req_1 : boolean;
  signal ptr_deref_1860_load_0_ack_1 : boolean;
  signal ptr_deref_1933_load_0_req_0 : boolean;
  signal ptr_deref_1933_load_0_ack_0 : boolean;
  signal ptr_deref_1933_load_0_req_1 : boolean;
  signal ptr_deref_1933_load_0_ack_1 : boolean;
  signal ptr_deref_1945_load_0_req_0 : boolean;
  signal ptr_deref_1945_load_0_ack_0 : boolean;
  signal ptr_deref_1945_load_0_req_1 : boolean;
  signal ptr_deref_1945_load_0_ack_1 : boolean;
  signal type_cast_1972_inst_req_0 : boolean;
  signal type_cast_1972_inst_ack_0 : boolean;
  signal type_cast_1972_inst_req_1 : boolean;
  signal type_cast_1972_inst_ack_1 : boolean;
  signal type_cast_1977_inst_req_0 : boolean;
  signal type_cast_1977_inst_ack_0 : boolean;
  signal type_cast_1977_inst_req_1 : boolean;
  signal type_cast_1977_inst_ack_1 : boolean;
  signal type_cast_2099_inst_req_0 : boolean;
  signal type_cast_2099_inst_ack_0 : boolean;
  signal type_cast_2099_inst_req_1 : boolean;
  signal type_cast_2099_inst_ack_1 : boolean;
  signal type_cast_2129_inst_req_0 : boolean;
  signal type_cast_2129_inst_ack_0 : boolean;
  signal type_cast_2129_inst_req_1 : boolean;
  signal type_cast_2129_inst_ack_1 : boolean;
  signal array_obj_ref_2135_index_offset_req_0 : boolean;
  signal array_obj_ref_2135_index_offset_ack_0 : boolean;
  signal array_obj_ref_2135_index_offset_req_1 : boolean;
  signal array_obj_ref_2135_index_offset_ack_1 : boolean;
  signal addr_of_2136_final_reg_req_0 : boolean;
  signal addr_of_2136_final_reg_ack_0 : boolean;
  signal addr_of_2136_final_reg_req_1 : boolean;
  signal addr_of_2136_final_reg_ack_1 : boolean;
  signal ptr_deref_2140_load_0_req_0 : boolean;
  signal ptr_deref_2140_load_0_ack_0 : boolean;
  signal ptr_deref_2140_load_0_req_1 : boolean;
  signal ptr_deref_2140_load_0_ack_1 : boolean;
  signal type_cast_2160_inst_req_0 : boolean;
  signal type_cast_2160_inst_ack_0 : boolean;
  signal type_cast_2160_inst_req_1 : boolean;
  signal type_cast_2160_inst_ack_1 : boolean;
  signal array_obj_ref_2166_index_offset_req_0 : boolean;
  signal array_obj_ref_2166_index_offset_ack_0 : boolean;
  signal array_obj_ref_2166_index_offset_req_1 : boolean;
  signal array_obj_ref_2166_index_offset_ack_1 : boolean;
  signal addr_of_2167_final_reg_req_0 : boolean;
  signal addr_of_2167_final_reg_ack_0 : boolean;
  signal addr_of_2167_final_reg_req_1 : boolean;
  signal addr_of_2167_final_reg_ack_1 : boolean;
  signal ptr_deref_2170_store_0_req_0 : boolean;
  signal ptr_deref_2170_store_0_ack_0 : boolean;
  signal ptr_deref_2170_store_0_req_1 : boolean;
  signal ptr_deref_2170_store_0_ack_1 : boolean;
  signal type_cast_2176_inst_req_0 : boolean;
  signal type_cast_2176_inst_ack_0 : boolean;
  signal type_cast_2176_inst_req_1 : boolean;
  signal type_cast_2176_inst_ack_1 : boolean;
  signal if_stmt_2189_branch_req_0 : boolean;
  signal if_stmt_2189_branch_ack_1 : boolean;
  signal if_stmt_2189_branch_ack_0 : boolean;
  signal type_cast_2213_inst_req_0 : boolean;
  signal type_cast_2213_inst_ack_0 : boolean;
  signal type_cast_2213_inst_req_1 : boolean;
  signal type_cast_2213_inst_ack_1 : boolean;
  signal if_stmt_2220_branch_req_0 : boolean;
  signal if_stmt_2220_branch_ack_1 : boolean;
  signal if_stmt_2220_branch_ack_0 : boolean;
  signal type_cast_2241_inst_req_0 : boolean;
  signal type_cast_2241_inst_ack_0 : boolean;
  signal type_cast_2241_inst_req_1 : boolean;
  signal type_cast_2241_inst_ack_1 : boolean;
  signal type_cast_2261_inst_req_0 : boolean;
  signal type_cast_2261_inst_ack_0 : boolean;
  signal type_cast_2261_inst_req_1 : boolean;
  signal type_cast_2261_inst_ack_1 : boolean;
  signal if_stmt_2268_branch_req_0 : boolean;
  signal if_stmt_2268_branch_ack_1 : boolean;
  signal if_stmt_2268_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2276_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2276_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2276_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2276_inst_ack_1 : boolean;
  signal phi_stmt_1961_req_1 : boolean;
  signal type_cast_1958_inst_req_0 : boolean;
  signal type_cast_1958_inst_ack_0 : boolean;
  signal type_cast_1958_inst_req_1 : boolean;
  signal type_cast_1958_inst_ack_1 : boolean;
  signal phi_stmt_1955_req_0 : boolean;
  signal type_cast_1964_inst_req_0 : boolean;
  signal type_cast_1964_inst_ack_0 : boolean;
  signal type_cast_1964_inst_req_1 : boolean;
  signal type_cast_1964_inst_ack_1 : boolean;
  signal phi_stmt_1961_req_0 : boolean;
  signal type_cast_1960_inst_req_0 : boolean;
  signal type_cast_1960_inst_ack_0 : boolean;
  signal type_cast_1960_inst_req_1 : boolean;
  signal type_cast_1960_inst_ack_1 : boolean;
  signal phi_stmt_1955_req_1 : boolean;
  signal phi_stmt_1955_ack_0 : boolean;
  signal phi_stmt_1961_ack_0 : boolean;
  signal type_cast_2086_inst_req_0 : boolean;
  signal type_cast_2086_inst_ack_0 : boolean;
  signal type_cast_2086_inst_req_1 : boolean;
  signal type_cast_2086_inst_ack_1 : boolean;
  signal phi_stmt_2083_req_0 : boolean;
  signal phi_stmt_2083_req_1 : boolean;
  signal phi_stmt_2083_ack_0 : boolean;
  signal type_cast_2248_inst_req_0 : boolean;
  signal type_cast_2248_inst_ack_0 : boolean;
  signal type_cast_2248_inst_req_1 : boolean;
  signal type_cast_2248_inst_ack_1 : boolean;
  signal phi_stmt_2245_req_0 : boolean;
  signal type_cast_2256_inst_req_0 : boolean;
  signal type_cast_2256_inst_ack_0 : boolean;
  signal type_cast_2256_inst_req_1 : boolean;
  signal type_cast_2256_inst_ack_1 : boolean;
  signal phi_stmt_2251_req_1 : boolean;
  signal type_cast_2250_inst_req_0 : boolean;
  signal type_cast_2250_inst_ack_0 : boolean;
  signal type_cast_2250_inst_req_1 : boolean;
  signal type_cast_2250_inst_ack_1 : boolean;
  signal phi_stmt_2245_req_1 : boolean;
  signal type_cast_2254_inst_req_0 : boolean;
  signal type_cast_2254_inst_ack_0 : boolean;
  signal type_cast_2254_inst_req_1 : boolean;
  signal type_cast_2254_inst_ack_1 : boolean;
  signal phi_stmt_2251_req_0 : boolean;
  signal phi_stmt_2245_ack_0 : boolean;
  signal phi_stmt_2251_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_5207_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_5207_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_5207_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_5207_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_5207: Block -- control-path 
    signal convTransposeB_CP_5207_elements: BooleanArray(112 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_5207_elements(0) <= convTransposeB_CP_5207_start;
    convTransposeB_CP_5207_symbol <= convTransposeB_CP_5207_elements(72);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1813/$entry
      -- CP-element group 0: 	 branch_block_stmt_1813/branch_block_stmt_1813__entry__
      -- CP-element group 0: 	 branch_block_stmt_1813/assign_stmt_1816__entry__
      -- CP-element group 0: 	 branch_block_stmt_1813/assign_stmt_1816/$entry
      -- CP-element group 0: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_Sample/rr
      -- 
    rr_5265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(0), ack => RPIPE_Block1_start_1815_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_Update/cr
      -- 
    ra_5266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1815_inst_ack_0, ack => convTransposeB_CP_5207_elements(1)); -- 
    cr_5270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(1), ack => RPIPE_Block1_start_1815_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2:  members (265) 
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1816__exit__
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952__entry__
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1816/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1816/RPIPE_Block1_start_1815_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/word_access_complete/word_0/cr
      -- 
    ca_5271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1815_inst_ack_1, ack => convTransposeB_CP_5207_elements(2)); -- 
    cr_5548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => type_cast_1883_inst_req_1); -- 
    rr_5646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1909_load_0_req_0); -- 
    cr_5529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => LOAD_padding_1879_load_0_req_1); -- 
    cr_5657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1909_load_0_req_1); -- 
    cr_5612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => type_cast_1897_inst_req_1); -- 
    cr_5593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1893_load_0_req_1); -- 
    cr_5451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => type_cast_1864_inst_req_1); -- 
    cr_5496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1876_load_0_req_1); -- 
    rr_5518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => LOAD_padding_1879_load_0_req_0); -- 
    rr_5485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1876_load_0_req_0); -- 
    cr_5707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1921_load_0_req_1); -- 
    rr_5582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1893_load_0_req_0); -- 
    rr_5696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1921_load_0_req_0); -- 
    rr_5307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1828_load_0_req_0); -- 
    cr_5318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1828_load_0_req_1); -- 
    cr_5337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => type_cast_1838_inst_req_1); -- 
    rr_5371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1850_load_0_req_0); -- 
    cr_5382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1850_load_0_req_1); -- 
    rr_5421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1860_load_0_req_0); -- 
    cr_5432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1860_load_0_req_1); -- 
    rr_5746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1933_load_0_req_0); -- 
    cr_5757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1933_load_0_req_1); -- 
    rr_5796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1945_load_0_req_0); -- 
    cr_5807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1945_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Sample/word_access_start/word_0/ra
      -- 
    ra_5308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1828_load_0_ack_0, ack => convTransposeB_CP_5207_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/ptr_deref_1828_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/ptr_deref_1828_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/ptr_deref_1828_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1828_Update/ptr_deref_1828_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_Sample/rr
      -- 
    ca_5319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1828_load_0_ack_1, ack => convTransposeB_CP_5207_elements(4)); -- 
    rr_5332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(4), ack => type_cast_1838_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_Sample/ra
      -- 
    ra_5333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1838_inst_ack_0, ack => convTransposeB_CP_5207_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1838_Update/ca
      -- 
    ca_5338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1838_inst_ack_1, ack => convTransposeB_CP_5207_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Sample/word_access_start/word_0/ra
      -- 
    ra_5372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1850_load_0_ack_0, ack => convTransposeB_CP_5207_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	31 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/ptr_deref_1850_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/ptr_deref_1850_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/ptr_deref_1850_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1850_Update/ptr_deref_1850_Merge/merge_ack
      -- 
    ca_5383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1850_load_0_ack_1, ack => convTransposeB_CP_5207_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Sample/word_access_start/word_0/ra
      -- 
    ra_5422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1860_load_0_ack_0, ack => convTransposeB_CP_5207_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (12) 
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/ptr_deref_1860_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/ptr_deref_1860_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/ptr_deref_1860_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1860_Update/ptr_deref_1860_Merge/merge_req
      -- 
    ca_5433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1860_load_0_ack_1, ack => convTransposeB_CP_5207_elements(10)); -- 
    rr_5446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(10), ack => type_cast_1864_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_sample_completed_
      -- 
    ra_5447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1864_inst_ack_0, ack => convTransposeB_CP_5207_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	31 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1864_Update/ca
      -- 
    ca_5452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1864_inst_ack_1, ack => convTransposeB_CP_5207_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_sample_completed_
      -- 
    ra_5486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1876_load_0_ack_0, ack => convTransposeB_CP_5207_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/ptr_deref_1876_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/ptr_deref_1876_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/ptr_deref_1876_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/ptr_deref_1876_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1876_update_completed_
      -- 
    ca_5497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1876_load_0_ack_1, ack => convTransposeB_CP_5207_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Sample/word_access_start/$exit
      -- 
    ra_5519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1879_load_0_ack_0, ack => convTransposeB_CP_5207_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (12) 
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/LOAD_padding_1879_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/LOAD_padding_1879_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/LOAD_padding_1879_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/LOAD_padding_1879_Merge/merge_ack
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/LOAD_padding_1879_update_completed_
      -- 
    ca_5530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1879_load_0_ack_1, ack => convTransposeB_CP_5207_elements(16)); -- 
    rr_5543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(16), ack => type_cast_1883_inst_req_0); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_sample_completed_
      -- 
    ra_5544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1883_inst_ack_0, ack => convTransposeB_CP_5207_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	31 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1883_Update/$exit
      -- 
    ca_5549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1883_inst_ack_1, ack => convTransposeB_CP_5207_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Sample/word_access_start/word_0/ra
      -- CP-element group 19: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Sample/word_access_start/word_0/$exit
      -- 
    ra_5583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1893_load_0_ack_0, ack => convTransposeB_CP_5207_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/ptr_deref_1893_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/ptr_deref_1893_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/ptr_deref_1893_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/ptr_deref_1893_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1893_Update/word_access_complete/word_0/$exit
      -- 
    ca_5594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1893_load_0_ack_1, ack => convTransposeB_CP_5207_elements(20)); -- 
    rr_5607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(20), ack => type_cast_1897_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_Sample/ra
      -- 
    ra_5608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1897_inst_ack_0, ack => convTransposeB_CP_5207_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	31 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/type_cast_1897_Update/ca
      -- 
    ca_5613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1897_inst_ack_1, ack => convTransposeB_CP_5207_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Sample/word_access_start/word_0/ra
      -- CP-element group 23: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Sample/word_access_start/$exit
      -- 
    ra_5647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1909_load_0_ack_0, ack => convTransposeB_CP_5207_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	31 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/ptr_deref_1909_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/ptr_deref_1909_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/ptr_deref_1909_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/ptr_deref_1909_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1909_Update/$exit
      -- 
    ca_5658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1909_load_0_ack_1, ack => convTransposeB_CP_5207_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Sample/word_access_start/word_0/ra
      -- CP-element group 25: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Sample/$exit
      -- 
    ra_5697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1921_load_0_ack_0, ack => convTransposeB_CP_5207_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/ptr_deref_1921_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/ptr_deref_1921_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/ptr_deref_1921_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1921_Update/ptr_deref_1921_Merge/merge_ack
      -- 
    ca_5708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1921_load_0_ack_1, ack => convTransposeB_CP_5207_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Sample/word_access_start/word_0/ra
      -- 
    ra_5747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1933_load_0_ack_0, ack => convTransposeB_CP_5207_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/ptr_deref_1933_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/ptr_deref_1933_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/ptr_deref_1933_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1933_Update/ptr_deref_1933_Merge/merge_ack
      -- 
    ca_5758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1933_load_0_ack_1, ack => convTransposeB_CP_5207_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Sample/word_access_start/word_0/ra
      -- 
    ra_5797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1945_load_0_ack_0, ack => convTransposeB_CP_5207_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/ptr_deref_1945_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/ptr_deref_1945_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/ptr_deref_1945_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/ptr_deref_1945_Update/ptr_deref_1945_Merge/merge_ack
      -- 
    ca_5808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1945_load_0_ack_1, ack => convTransposeB_CP_5207_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	12 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	18 
    -- CP-element group 31: 	24 
    -- CP-element group 31: 	22 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	6 
    -- CP-element group 31: 	8 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	73 
    -- CP-element group 31: 	74 
    -- CP-element group 31: 	75 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952__exit__
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1813/assign_stmt_1825_to_assign_stmt_1952/$exit
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/$entry
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/$entry
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/$entry
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/SplitProtocol/Update/cr
      -- 
    rr_6250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(31), ack => type_cast_1958_inst_req_0); -- 
    cr_6255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(31), ack => type_cast_1958_inst_req_1); -- 
    convTransposeB_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(12) & convTransposeB_CP_5207_elements(26) & convTransposeB_CP_5207_elements(18) & convTransposeB_CP_5207_elements(24) & convTransposeB_CP_5207_elements(22) & convTransposeB_CP_5207_elements(28) & convTransposeB_CP_5207_elements(30) & convTransposeB_CP_5207_elements(14) & convTransposeB_CP_5207_elements(6) & convTransposeB_CP_5207_elements(8);
      gj_convTransposeB_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	88 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_Sample/ra
      -- 
    ra_5825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1972_inst_ack_0, ack => convTransposeB_CP_5207_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	88 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_Update/ca
      -- 
    ca_5830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1972_inst_ack_1, ack => convTransposeB_CP_5207_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	88 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_Sample/ra
      -- 
    ra_5839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1977_inst_ack_0, ack => convTransposeB_CP_5207_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_Update/ca
      -- 
    ca_5844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1977_inst_ack_1, ack => convTransposeB_CP_5207_elements(35)); -- 
    -- CP-element group 36:  join  transition  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	92 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080__exit__
      -- CP-element group 36: 	 branch_block_stmt_1813/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 36: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/$exit
      -- CP-element group 36: 	 branch_block_stmt_1813/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_1813/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2083/$entry
      -- CP-element group 36: 	 branch_block_stmt_1813/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/$entry
      -- 
    convTransposeB_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(33) & convTransposeB_CP_5207_elements(35);
      gj_convTransposeB_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	94 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_Sample/ra
      -- 
    ra_5856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2099_inst_ack_0, ack => convTransposeB_CP_5207_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	94 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	47 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_Sample/rr
      -- 
    ca_5861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2099_inst_ack_1, ack => convTransposeB_CP_5207_elements(38)); -- 
    rr_5979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(38), ack => type_cast_2160_inst_req_0); -- 
    rr_5869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(38), ack => type_cast_2129_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_Sample/ra
      -- 
    ra_5870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2129_inst_ack_0, ack => convTransposeB_CP_5207_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	94 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (16) 
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_resized_1
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_scaled_1
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_computed_1
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_resize_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_resize_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_resize_1/index_resize_req
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_resize_1/index_resize_ack
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_scale_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_scale_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_scale_1/scale_rename_req
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_index_scale_1/scale_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_final_index_sum_regn_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_final_index_sum_regn_Sample/req
      -- 
    ca_5875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2129_inst_ack_1, ack => convTransposeB_CP_5207_elements(40)); -- 
    req_5900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(40), ack => array_obj_ref_2135_index_offset_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_final_index_sum_regn_sample_complete
      -- CP-element group 41: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_final_index_sum_regn_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_final_index_sum_regn_Sample/ack
      -- 
    ack_5901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2135_index_offset_ack_0, ack => convTransposeB_CP_5207_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	94 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_offset_calculated
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_final_index_sum_regn_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_final_index_sum_regn_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_request/$entry
      -- CP-element group 42: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_request/req
      -- 
    ack_5906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2135_index_offset_ack_1, ack => convTransposeB_CP_5207_elements(42)); -- 
    req_5915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(42), ack => addr_of_2136_final_reg_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_request/$exit
      -- CP-element group 43: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_request/ack
      -- 
    ack_5916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2136_final_reg_ack_0, ack => convTransposeB_CP_5207_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	94 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (24) 
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_complete/ack
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_base_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_word_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_base_address_resized
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_base_addr_resize/$entry
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_base_addr_resize/$exit
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_base_addr_resize/base_resize_req
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_base_addr_resize/base_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_word_addrgen/$entry
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_word_addrgen/$exit
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_word_addrgen/root_register_req
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_word_addrgen/root_register_ack
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Sample/word_access_start/word_0/rr
      -- 
    ack_5921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2136_final_reg_ack_1, ack => convTransposeB_CP_5207_elements(44)); -- 
    rr_5954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(44), ack => ptr_deref_2140_load_0_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Sample/word_access_start/word_0/ra
      -- 
    ra_5955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2140_load_0_ack_0, ack => convTransposeB_CP_5207_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	94 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	53 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/ptr_deref_2140_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/ptr_deref_2140_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/ptr_deref_2140_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/ptr_deref_2140_Merge/merge_ack
      -- 
    ca_5966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2140_load_0_ack_1, ack => convTransposeB_CP_5207_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_Sample/ra
      -- 
    ra_5980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2160_inst_ack_0, ack => convTransposeB_CP_5207_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	94 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (16) 
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_resized_1
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_scaled_1
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_computed_1
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_resize_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_resize_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_resize_1/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_resize_1/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_scale_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_scale_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_scale_1/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_index_scale_1/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_final_index_sum_regn_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_final_index_sum_regn_Sample/req
      -- 
    ca_5985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2160_inst_ack_1, ack => convTransposeB_CP_5207_elements(48)); -- 
    req_6010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(48), ack => array_obj_ref_2166_index_offset_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_final_index_sum_regn_sample_complete
      -- CP-element group 49: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_final_index_sum_regn_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_final_index_sum_regn_Sample/ack
      -- 
    ack_6011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2166_index_offset_ack_0, ack => convTransposeB_CP_5207_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	94 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (11) 
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_offset_calculated
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_final_index_sum_regn_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_final_index_sum_regn_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_request/$entry
      -- CP-element group 50: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_request/req
      -- 
    ack_6016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2166_index_offset_ack_1, ack => convTransposeB_CP_5207_elements(50)); -- 
    req_6025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(50), ack => addr_of_2167_final_reg_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_request/$exit
      -- CP-element group 51: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_request/ack
      -- 
    ack_6026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2167_final_reg_ack_0, ack => convTransposeB_CP_5207_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	94 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (19) 
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_complete/ack
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_word_addrgen/root_register_ack
      -- 
    ack_6031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2167_final_reg_ack_1, ack => convTransposeB_CP_5207_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	46 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/ptr_deref_2170_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/ptr_deref_2170_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/ptr_deref_2170_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/ptr_deref_2170_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/word_access_start/word_0/rr
      -- 
    rr_6069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(53), ack => ptr_deref_2170_store_0_req_0); -- 
    convTransposeB_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(46) & convTransposeB_CP_5207_elements(52);
      gj_convTransposeB_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Sample/word_access_start/word_0/ra
      -- 
    ra_6070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2170_store_0_ack_0, ack => convTransposeB_CP_5207_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	94 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Update/word_access_complete/word_0/ca
      -- 
    ca_6081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2170_store_0_ack_1, ack => convTransposeB_CP_5207_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	94 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_Sample/ra
      -- 
    ra_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2176_inst_ack_0, ack => convTransposeB_CP_5207_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	94 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_Update/ca
      -- 
    ca_6095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2176_inst_ack_1, ack => convTransposeB_CP_5207_elements(57)); -- 
    -- CP-element group 58:  branch  join  transition  place  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188__exit__
      -- CP-element group 58: 	 branch_block_stmt_1813/if_stmt_2189__entry__
      -- CP-element group 58: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/$exit
      -- CP-element group 58: 	 branch_block_stmt_1813/if_stmt_2189_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1813/if_stmt_2189_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_1813/if_stmt_2189_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_1813/if_stmt_2189_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_1813/R_cmp_2190_place
      -- CP-element group 58: 	 branch_block_stmt_1813/if_stmt_2189_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1813/if_stmt_2189_else_link/$entry
      -- 
    branch_req_6103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(58), ack => if_stmt_2189_branch_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(41) & convTransposeB_CP_5207_elements(55) & convTransposeB_CP_5207_elements(49) & convTransposeB_CP_5207_elements(57);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	89 
    -- CP-element group 59: 	90 
    -- CP-element group 59:  members (24) 
      -- CP-element group 59: 	 branch_block_stmt_1813/merge_stmt_2195__exit__
      -- CP-element group 59: 	 branch_block_stmt_1813/assign_stmt_2201__entry__
      -- CP-element group 59: 	 branch_block_stmt_1813/assign_stmt_2201__exit__
      -- CP-element group 59: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody
      -- CP-element group 59: 	 branch_block_stmt_1813/if_stmt_2189_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1813/if_stmt_2189_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1813/whilex_xbody_ifx_xthen
      -- CP-element group 59: 	 branch_block_stmt_1813/assign_stmt_2201/$entry
      -- CP-element group 59: 	 branch_block_stmt_1813/assign_stmt_2201/$exit
      -- CP-element group 59: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/$entry
      -- CP-element group 59: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/$entry
      -- CP-element group 59: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_1813/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1813/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1813/merge_stmt_2195_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1813/merge_stmt_2195_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1813/merge_stmt_2195_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1813/merge_stmt_2195_PhiAck/dummy
      -- 
    if_choice_transition_6108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2189_branch_ack_1, ack => convTransposeB_CP_5207_elements(59)); -- 
    rr_6331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(59), ack => type_cast_2086_inst_req_0); -- 
    cr_6336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(59), ack => type_cast_2086_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (18) 
      -- CP-element group 60: 	 branch_block_stmt_1813/merge_stmt_2203__exit__
      -- CP-element group 60: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219__entry__
      -- CP-element group 60: 	 branch_block_stmt_1813/if_stmt_2189_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_1813/if_stmt_2189_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_1813/whilex_xbody_ifx_xelse
      -- CP-element group 60: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/$entry
      -- CP-element group 60: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_1813/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_1813/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_1813/merge_stmt_2203_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_1813/merge_stmt_2203_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_1813/merge_stmt_2203_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_1813/merge_stmt_2203_PhiAck/dummy
      -- 
    else_choice_transition_6112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2189_branch_ack_0, ack => convTransposeB_CP_5207_elements(60)); -- 
    rr_6128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(60), ack => type_cast_2213_inst_req_0); -- 
    cr_6133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(60), ack => type_cast_2213_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_Sample/ra
      -- 
    ra_6129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2213_inst_ack_0, ack => convTransposeB_CP_5207_elements(61)); -- 
    -- CP-element group 62:  branch  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (13) 
      -- CP-element group 62: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219__exit__
      -- CP-element group 62: 	 branch_block_stmt_1813/if_stmt_2220__entry__
      -- CP-element group 62: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/$exit
      -- CP-element group 62: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1813/assign_stmt_2209_to_assign_stmt_2219/type_cast_2213_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1813/if_stmt_2220_dead_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1813/if_stmt_2220_eval_test/$entry
      -- CP-element group 62: 	 branch_block_stmt_1813/if_stmt_2220_eval_test/$exit
      -- CP-element group 62: 	 branch_block_stmt_1813/if_stmt_2220_eval_test/branch_req
      -- CP-element group 62: 	 branch_block_stmt_1813/R_cmp77_2221_place
      -- CP-element group 62: 	 branch_block_stmt_1813/if_stmt_2220_if_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1813/if_stmt_2220_else_link/$entry
      -- 
    ca_6134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2213_inst_ack_1, ack => convTransposeB_CP_5207_elements(62)); -- 
    branch_req_6142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(62), ack => if_stmt_2220_branch_req_0); -- 
    -- CP-element group 63:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (18) 
      -- CP-element group 63: 	 branch_block_stmt_1813/merge_stmt_2226__exit__
      -- CP-element group 63: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242__entry__
      -- CP-element group 63: 	 branch_block_stmt_1813/if_stmt_2220_if_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_1813/if_stmt_2220_if_link/if_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_1813/ifx_xelse_ifx_xthen79
      -- CP-element group 63: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/$entry
      -- CP-element group 63: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_Update/cr
      -- CP-element group 63: 	 branch_block_stmt_1813/ifx_xelse_ifx_xthen79_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_1813/ifx_xelse_ifx_xthen79_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_1813/merge_stmt_2226_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_1813/merge_stmt_2226_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_1813/merge_stmt_2226_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_1813/merge_stmt_2226_PhiAck/dummy
      -- 
    if_choice_transition_6147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2220_branch_ack_1, ack => convTransposeB_CP_5207_elements(63)); -- 
    rr_6164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(63), ack => type_cast_2241_inst_req_0); -- 
    cr_6169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(63), ack => type_cast_2241_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	95 
    -- CP-element group 64: 	96 
    -- CP-element group 64: 	98 
    -- CP-element group 64: 	99 
    -- CP-element group 64:  members (20) 
      -- CP-element group 64: 	 branch_block_stmt_1813/if_stmt_2220_else_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1813/if_stmt_2220_else_link/else_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2220_branch_ack_0, ack => convTransposeB_CP_5207_elements(64)); -- 
    rr_6405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(64), ack => type_cast_2248_inst_req_0); -- 
    cr_6410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(64), ack => type_cast_2248_inst_req_1); -- 
    rr_6428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(64), ack => type_cast_2256_inst_req_0); -- 
    cr_6433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(64), ack => type_cast_2256_inst_req_1); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_Sample/ra
      -- 
    ra_6165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2241_inst_ack_0, ack => convTransposeB_CP_5207_elements(65)); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	105 
    -- CP-element group 66: 	106 
    -- CP-element group 66: 	102 
    -- CP-element group 66: 	103 
    -- CP-element group 66:  members (23) 
      -- CP-element group 66: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242__exit__
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend
      -- CP-element group 66: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/$exit
      -- CP-element group 66: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1813/assign_stmt_2232_to_assign_stmt_2242/type_cast_2241_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Update/cr
      -- 
    ca_6170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2241_inst_ack_1, ack => convTransposeB_CP_5207_elements(66)); -- 
    rr_6454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(66), ack => type_cast_2250_inst_req_0); -- 
    cr_6459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(66), ack => type_cast_2250_inst_req_1); -- 
    rr_6477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(66), ack => type_cast_2254_inst_req_0); -- 
    cr_6482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(66), ack => type_cast_2254_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	112 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_Sample/ra
      -- 
    ra_6182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2261_inst_ack_0, ack => convTransposeB_CP_5207_elements(67)); -- 
    -- CP-element group 68:  branch  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	112 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (13) 
      -- CP-element group 68: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267__exit__
      -- CP-element group 68: 	 branch_block_stmt_1813/if_stmt_2268__entry__
      -- CP-element group 68: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/$exit
      -- CP-element group 68: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_1813/if_stmt_2268_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1813/if_stmt_2268_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1813/if_stmt_2268_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1813/if_stmt_2268_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1813/R_cmp89_2269_place
      -- CP-element group 68: 	 branch_block_stmt_1813/if_stmt_2268_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1813/if_stmt_2268_else_link/$entry
      -- 
    ca_6187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2261_inst_ack_1, ack => convTransposeB_CP_5207_elements(68)); -- 
    branch_req_6195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(68), ack => if_stmt_2268_branch_req_0); -- 
    -- CP-element group 69:  merge  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (15) 
      -- CP-element group 69: 	 branch_block_stmt_1813/merge_stmt_2274__exit__
      -- CP-element group 69: 	 branch_block_stmt_1813/assign_stmt_2278__entry__
      -- CP-element group 69: 	 branch_block_stmt_1813/if_stmt_2268_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1813/if_stmt_2268_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1813/ifx_xend_whilex_xend
      -- CP-element group 69: 	 branch_block_stmt_1813/assign_stmt_2278/$entry
      -- CP-element group 69: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_Sample/req
      -- CP-element group 69: 	 branch_block_stmt_1813/ifx_xend_whilex_xend_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1813/ifx_xend_whilex_xend_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1813/merge_stmt_2274_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1813/merge_stmt_2274_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1813/merge_stmt_2274_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1813/merge_stmt_2274_PhiAck/dummy
      -- 
    if_choice_transition_6200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2268_branch_ack_1, ack => convTransposeB_CP_5207_elements(69)); -- 
    req_6217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(69), ack => WPIPE_Block1_done_2276_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	81 
    -- CP-element group 70: 	82 
    -- CP-element group 70: 	78 
    -- CP-element group 70: 	79 
    -- CP-element group 70:  members (20) 
      -- CP-element group 70: 	 branch_block_stmt_1813/if_stmt_2268_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1813/if_stmt_2268_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/SplitProtocol/Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2268_branch_ack_0, ack => convTransposeB_CP_5207_elements(70)); -- 
    rr_6276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(70), ack => type_cast_1964_inst_req_0); -- 
    cr_6281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(70), ack => type_cast_1964_inst_req_1); -- 
    rr_6299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(70), ack => type_cast_1960_inst_req_0); -- 
    cr_6304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(70), ack => type_cast_1960_inst_req_1); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_Sample/ack
      -- CP-element group 71: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_Update/req
      -- 
    ack_6218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2276_inst_ack_0, ack => convTransposeB_CP_5207_elements(71)); -- 
    req_6222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(71), ack => WPIPE_Block1_done_2276_inst_req_1); -- 
    -- CP-element group 72:  transition  place  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (16) 
      -- CP-element group 72: 	 $exit
      -- CP-element group 72: 	 branch_block_stmt_1813/$exit
      -- CP-element group 72: 	 branch_block_stmt_1813/branch_block_stmt_1813__exit__
      -- CP-element group 72: 	 branch_block_stmt_1813/assign_stmt_2278__exit__
      -- CP-element group 72: 	 branch_block_stmt_1813/return__
      -- CP-element group 72: 	 branch_block_stmt_1813/merge_stmt_2280__exit__
      -- CP-element group 72: 	 branch_block_stmt_1813/assign_stmt_2278/$exit
      -- CP-element group 72: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1813/assign_stmt_2278/WPIPE_Block1_done_2276_Update/ack
      -- CP-element group 72: 	 branch_block_stmt_1813/return___PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_1813/return___PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_1813/merge_stmt_2280_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1813/merge_stmt_2280_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_1813/merge_stmt_2280_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_1813/merge_stmt_2280_PhiAck/dummy
      -- 
    ack_6223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2276_inst_ack_1, ack => convTransposeB_CP_5207_elements(72)); -- 
    -- CP-element group 73:  transition  output  delay-element  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	31 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/$exit
      -- CP-element group 73: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1967_konst_delay_trans
      -- CP-element group 73: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_req
      -- 
    phi_stmt_1961_req_6234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1961_req_6234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(73), ack => phi_stmt_1961_req_1); -- 
    -- Element group convTransposeB_CP_5207_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => convTransposeB_CP_5207_elements(31), ack => convTransposeB_CP_5207_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	31 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/SplitProtocol/Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/SplitProtocol/Sample/ra
      -- 
    ra_6251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1958_inst_ack_0, ack => convTransposeB_CP_5207_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	31 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/SplitProtocol/Update/ca
      -- 
    ca_6256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1958_inst_ack_1, ack => convTransposeB_CP_5207_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/$exit
      -- CP-element group 76: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/$exit
      -- CP-element group 76: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1958/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_req
      -- 
    phi_stmt_1955_req_6257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1955_req_6257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(76), ack => phi_stmt_1955_req_0); -- 
    convTransposeB_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(74) & convTransposeB_CP_5207_elements(75);
      gj_convTransposeB_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: 	73 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	85 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1813/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(76) & convTransposeB_CP_5207_elements(73);
      gj_convTransposeB_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	70 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/SplitProtocol/Sample/ra
      -- 
    ra_6277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1964_inst_ack_0, ack => convTransposeB_CP_5207_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	70 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/SplitProtocol/Update/ca
      -- 
    ca_6282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1964_inst_ack_1, ack => convTransposeB_CP_5207_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	84 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/$exit
      -- CP-element group 80: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/$exit
      -- CP-element group 80: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_sources/type_cast_1964/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1961/phi_stmt_1961_req
      -- 
    phi_stmt_1961_req_6283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1961_req_6283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(80), ack => phi_stmt_1961_req_0); -- 
    convTransposeB_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(78) & convTransposeB_CP_5207_elements(79);
      gj_convTransposeB_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	70 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/SplitProtocol/Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/SplitProtocol/Sample/ra
      -- 
    ra_6300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1960_inst_ack_0, ack => convTransposeB_CP_5207_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/SplitProtocol/Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/SplitProtocol/Update/ca
      -- 
    ca_6305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1960_inst_ack_1, ack => convTransposeB_CP_5207_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/$exit
      -- CP-element group 83: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/$exit
      -- CP-element group 83: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_sources/type_cast_1960/SplitProtocol/$exit
      -- CP-element group 83: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1955/phi_stmt_1955_req
      -- 
    phi_stmt_1955_req_6306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1955_req_6306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(83), ack => phi_stmt_1955_req_1); -- 
    convTransposeB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(81) & convTransposeB_CP_5207_elements(82);
      gj_convTransposeB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: 	80 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1813/ifx_xend_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(83) & convTransposeB_CP_5207_elements(80);
      gj_convTransposeB_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  merge  fork  transition  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	77 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1813/merge_stmt_1954_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_1813/merge_stmt_1954_PhiAck/$entry
      -- 
    convTransposeB_CP_5207_elements(85) <= OrReduce(convTransposeB_CP_5207_elements(77) & convTransposeB_CP_5207_elements(84));
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1813/merge_stmt_1954_PhiAck/phi_stmt_1955_ack
      -- 
    phi_stmt_1955_ack_6311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1955_ack_0, ack => convTransposeB_CP_5207_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1813/merge_stmt_1954_PhiAck/phi_stmt_1961_ack
      -- 
    phi_stmt_1961_ack_6312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1961_ack_0, ack => convTransposeB_CP_5207_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  place  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	32 
    -- CP-element group 88: 	33 
    -- CP-element group 88: 	34 
    -- CP-element group 88: 	35 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 branch_block_stmt_1813/merge_stmt_1954__exit__
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080__entry__
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/$entry
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1972_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1813/assign_stmt_1973_to_assign_stmt_2080/type_cast_1977_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1813/merge_stmt_1954_PhiAck/$exit
      -- 
    rr_5824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(88), ack => type_cast_1972_inst_req_0); -- 
    cr_5829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(88), ack => type_cast_1972_inst_req_1); -- 
    rr_5838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(88), ack => type_cast_1977_inst_req_0); -- 
    cr_5843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(88), ack => type_cast_1977_inst_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(86) & convTransposeB_CP_5207_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	59 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Sample/ra
      -- 
    ra_6332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2086_inst_ack_0, ack => convTransposeB_CP_5207_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	59 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/Update/ca
      -- 
    ca_6337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2086_inst_ack_1, ack => convTransposeB_CP_5207_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 91: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/$exit
      -- CP-element group 91: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/$exit
      -- CP-element group 91: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2086/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1813/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_req
      -- 
    phi_stmt_2083_req_6338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2083_req_6338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(91), ack => phi_stmt_2083_req_0); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(89) & convTransposeB_CP_5207_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  output  delay-element  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	36 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1813/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 92: 	 branch_block_stmt_1813/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2083/$exit
      -- CP-element group 92: 	 branch_block_stmt_1813/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1813/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_sources/type_cast_2089_konst_delay_trans
      -- CP-element group 92: 	 branch_block_stmt_1813/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2083/phi_stmt_2083_req
      -- 
    phi_stmt_2083_req_6349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2083_req_6349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(92), ack => phi_stmt_2083_req_1); -- 
    -- Element group convTransposeB_CP_5207_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => convTransposeB_CP_5207_elements(36), ack => convTransposeB_CP_5207_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  merge  transition  place  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1813/merge_stmt_2082_PhiReqMerge
      -- CP-element group 93: 	 branch_block_stmt_1813/merge_stmt_2082_PhiAck/$entry
      -- 
    convTransposeB_CP_5207_elements(93) <= OrReduce(convTransposeB_CP_5207_elements(92) & convTransposeB_CP_5207_elements(91));
    -- CP-element group 94:  fork  transition  place  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	42 
    -- CP-element group 94: 	44 
    -- CP-element group 94: 	48 
    -- CP-element group 94: 	40 
    -- CP-element group 94: 	46 
    -- CP-element group 94: 	52 
    -- CP-element group 94: 	55 
    -- CP-element group 94: 	50 
    -- CP-element group 94: 	56 
    -- CP-element group 94: 	57 
    -- CP-element group 94: 	37 
    -- CP-element group 94: 	38 
    -- CP-element group 94:  members (45) 
      -- CP-element group 94: 	 branch_block_stmt_1813/merge_stmt_2082__exit__
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188__entry__
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2099_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2129_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_final_index_sum_regn_update_start
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_final_index_sum_regn_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2135_final_index_sum_regn_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2136_complete/req
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2140_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2160_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_final_index_sum_regn_update_start
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_final_index_sum_regn_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/array_obj_ref_2166_final_index_sum_regn_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/addr_of_2167_complete/req
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/ptr_deref_2170_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1813/assign_stmt_2096_to_assign_stmt_2188/type_cast_2176_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1813/merge_stmt_2082_PhiAck/$exit
      -- CP-element group 94: 	 branch_block_stmt_1813/merge_stmt_2082_PhiAck/phi_stmt_2083_ack
      -- 
    phi_stmt_2083_ack_6354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2083_ack_0, ack => convTransposeB_CP_5207_elements(94)); -- 
    rr_5855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2099_inst_req_0); -- 
    cr_5860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2099_inst_req_1); -- 
    cr_5874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2129_inst_req_1); -- 
    req_5905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => array_obj_ref_2135_index_offset_req_1); -- 
    req_5920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => addr_of_2136_final_reg_req_1); -- 
    cr_5965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => ptr_deref_2140_load_0_req_1); -- 
    cr_5984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2160_inst_req_1); -- 
    req_6015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => array_obj_ref_2166_index_offset_req_1); -- 
    req_6030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => addr_of_2167_final_reg_req_1); -- 
    cr_6080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => ptr_deref_2170_store_0_req_1); -- 
    rr_6089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2176_inst_req_0); -- 
    cr_6094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2176_inst_req_1); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	64 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Sample/ra
      -- 
    ra_6406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2248_inst_ack_0, ack => convTransposeB_CP_5207_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	64 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/Update/ca
      -- 
    ca_6411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2248_inst_ack_1, ack => convTransposeB_CP_5207_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/$exit
      -- CP-element group 97: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/$exit
      -- CP-element group 97: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2248/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_req
      -- 
    phi_stmt_2245_req_6412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2245_req_6412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(97), ack => phi_stmt_2245_req_0); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(95) & convTransposeB_CP_5207_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	64 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/SplitProtocol/Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/SplitProtocol/Sample/ra
      -- 
    ra_6429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2256_inst_ack_0, ack => convTransposeB_CP_5207_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	64 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/SplitProtocol/Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/SplitProtocol/Update/ca
      -- 
    ca_6434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2256_inst_ack_1, ack => convTransposeB_CP_5207_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/$exit
      -- CP-element group 100: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/$exit
      -- CP-element group 100: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2256/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_req
      -- 
    phi_stmt_2251_req_6435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2251_req_6435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(100), ack => phi_stmt_2251_req_1); -- 
    convTransposeB_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(98) & convTransposeB_CP_5207_elements(99);
      gj_convTransposeB_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	109 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1813/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(97) & convTransposeB_CP_5207_elements(100);
      gj_convTransposeB_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	66 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Sample/ra
      -- 
    ra_6455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2250_inst_ack_0, ack => convTransposeB_CP_5207_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/Update/ca
      -- 
    ca_6460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2250_inst_ack_1, ack => convTransposeB_CP_5207_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/$exit
      -- CP-element group 104: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/$exit
      -- CP-element group 104: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_sources/type_cast_2250/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2245/phi_stmt_2245_req
      -- 
    phi_stmt_2245_req_6461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2245_req_6461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(104), ack => phi_stmt_2245_req_1); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(102) & convTransposeB_CP_5207_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	66 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Sample/ra
      -- 
    ra_6478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2254_inst_ack_0, ack => convTransposeB_CP_5207_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	66 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Update/ca
      -- 
    ca_6483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2254_inst_ack_1, ack => convTransposeB_CP_5207_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/$exit
      -- CP-element group 107: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/$exit
      -- CP-element group 107: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2251/phi_stmt_2251_req
      -- 
    phi_stmt_2251_req_6484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2251_req_6484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(107), ack => phi_stmt_2251_req_0); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(105) & convTransposeB_CP_5207_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: 	104 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1813/ifx_xthen79_ifx_xend_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(107) & convTransposeB_CP_5207_elements(104);
      gj_convTransposeB_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  merge  fork  transition  place  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: 	101 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1813/merge_stmt_2244_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_1813/merge_stmt_2244_PhiAck/$entry
      -- 
    convTransposeB_CP_5207_elements(109) <= OrReduce(convTransposeB_CP_5207_elements(108) & convTransposeB_CP_5207_elements(101));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1813/merge_stmt_2244_PhiAck/phi_stmt_2245_ack
      -- 
    phi_stmt_2245_ack_6489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2245_ack_0, ack => convTransposeB_CP_5207_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1813/merge_stmt_2244_PhiAck/phi_stmt_2251_ack
      -- 
    phi_stmt_2251_ack_6490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2251_ack_0, ack => convTransposeB_CP_5207_elements(111)); -- 
    -- CP-element group 112:  join  fork  transition  place  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: 	68 
    -- CP-element group 112:  members (10) 
      -- CP-element group 112: 	 branch_block_stmt_1813/merge_stmt_2244__exit__
      -- CP-element group 112: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267__entry__
      -- CP-element group 112: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/$entry
      -- CP-element group 112: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_update_start_
      -- CP-element group 112: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_1813/assign_stmt_2262_to_assign_stmt_2267/type_cast_2261_Update/cr
      -- CP-element group 112: 	 branch_block_stmt_1813/merge_stmt_2244_PhiAck/$exit
      -- 
    rr_6181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(112), ack => type_cast_2261_inst_req_0); -- 
    cr_6186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(112), ack => type_cast_2261_inst_req_1); -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(110) & convTransposeB_CP_5207_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(112), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2042_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2063_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2123_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2154_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1879_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1879_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom61_2165_resized : std_logic_vector(13 downto 0);
    signal R_idxprom61_2165_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2134_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2134_scaled : std_logic_vector(13 downto 0);
    signal add17_2105 : std_logic_vector(31 downto 0);
    signal add25_2003 : std_logic_vector(31 downto 0);
    signal add36_2018 : std_logic_vector(31 downto 0);
    signal add51_2075 : std_logic_vector(31 downto 0);
    signal add53_2110 : std_logic_vector(31 downto 0);
    signal add66_2183 : std_logic_vector(31 downto 0);
    signal add_1988 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2135_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2135_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2135_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2135_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2135_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2135_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2166_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2166_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2166_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2166_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2166_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2166_root_address : std_logic_vector(13 downto 0);
    signal arrayidx62_2168 : std_logic_vector(31 downto 0);
    signal arrayidx_2137 : std_logic_vector(31 downto 0);
    signal call_1816 : std_logic_vector(15 downto 0);
    signal cmp77_2219 : std_logic_vector(0 downto 0);
    signal cmp89_2267 : std_logic_vector(0 downto 0);
    signal cmp_2188 : std_logic_vector(0 downto 0);
    signal conv12_1973 : std_logic_vector(31 downto 0);
    signal conv15_1978 : std_logic_vector(31 downto 0);
    signal conv22_1865 : std_logic_vector(31 downto 0);
    signal conv27_1884 : std_logic_vector(31 downto 0);
    signal conv33_1898 : std_logic_vector(31 downto 0);
    signal conv46_2044 : std_logic_vector(31 downto 0);
    signal conv49_2065 : std_logic_vector(31 downto 0);
    signal conv65_2177 : std_logic_vector(31 downto 0);
    signal conv75_2214 : std_logic_vector(31 downto 0);
    signal conv84_2242 : std_logic_vector(15 downto 0);
    signal conv86_2262 : std_logic_vector(31 downto 0);
    signal conv9102_2100 : std_logic_vector(31 downto 0);
    signal conv_1839 : std_logic_vector(15 downto 0);
    signal div83_2238 : std_logic_vector(31 downto 0);
    signal div88_1952 : std_logic_vector(31 downto 0);
    signal div_1835 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1942 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1825 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1847 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1857 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1873 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1890 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1906 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1918 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1930 : std_logic_vector(31 downto 0);
    signal idxprom61_2161 : std_logic_vector(63 downto 0);
    signal idxprom_2130 : std_logic_vector(63 downto 0);
    signal inc81_2232 : std_logic_vector(15 downto 0);
    signal inc_2209 : std_logic_vector(15 downto 0);
    signal indvar_2083 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2201 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2251 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1961 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1955 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2245 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2096 : std_logic_vector(15 downto 0);
    signal mul16_1993 : std_logic_vector(31 downto 0);
    signal mul23_1998 : std_logic_vector(31 downto 0);
    signal mul34_2013 : std_logic_vector(31 downto 0);
    signal mul50_2070 : std_logic_vector(31 downto 0);
    signal mul52_2080 : std_logic_vector(31 downto 0);
    signal mul_1983 : std_logic_vector(31 downto 0);
    signal ptr_deref_1828_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1828_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1828_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1828_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1828_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1850_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1850_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1850_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1850_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1850_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1860_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1860_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1860_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1860_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1860_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1876_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1876_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1876_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1876_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1876_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1893_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1893_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1893_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1893_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1893_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1909_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1909_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1909_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1909_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1909_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1921_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1921_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1921_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1921_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1921_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1933_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1933_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1933_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1933_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1933_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1945_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1945_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1945_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1945_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1945_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2140_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2140_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2140_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2140_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2140_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2170_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2170_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2170_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2170_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2170_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2170_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext103_2056 : std_logic_vector(31 downto 0);
    signal sext105_2116 : std_logic_vector(31 downto 0);
    signal sext106_2147 : std_logic_vector(31 downto 0);
    signal sext_2035 : std_logic_vector(31 downto 0);
    signal shr60_2156 : std_logic_vector(31 downto 0);
    signal shr_2125 : std_logic_vector(31 downto 0);
    signal sub28_2050 : std_logic_vector(31 downto 0);
    signal sub39_2023 : std_logic_vector(31 downto 0);
    signal sub40_2029 : std_logic_vector(31 downto 0);
    signal sub_2008 : std_logic_vector(31 downto 0);
    signal tmp10_1851 : std_logic_vector(31 downto 0);
    signal tmp21_1861 : std_logic_vector(15 downto 0);
    signal tmp24_1877 : std_logic_vector(31 downto 0);
    signal tmp26_1880 : std_logic_vector(15 downto 0);
    signal tmp32_1894 : std_logic_vector(15 downto 0);
    signal tmp35_1910 : std_logic_vector(31 downto 0);
    signal tmp44_1922 : std_logic_vector(31 downto 0);
    signal tmp47_1934 : std_logic_vector(31 downto 0);
    signal tmp57_2141 : std_logic_vector(63 downto 0);
    signal tmp87_1946 : std_logic_vector(31 downto 0);
    signal tmp_1829 : std_logic_vector(31 downto 0);
    signal type_cast_1833_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1950_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1958_wire : std_logic_vector(15 downto 0);
    signal type_cast_1960_wire : std_logic_vector(15 downto 0);
    signal type_cast_1964_wire : std_logic_vector(15 downto 0);
    signal type_cast_1967_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1971_wire : std_logic_vector(31 downto 0);
    signal type_cast_1976_wire : std_logic_vector(31 downto 0);
    signal type_cast_2027_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2033_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2038_wire : std_logic_vector(31 downto 0);
    signal type_cast_2041_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2048_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2054_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2059_wire : std_logic_vector(31 downto 0);
    signal type_cast_2062_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2086_wire : std_logic_vector(15 downto 0);
    signal type_cast_2089_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2094_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2114_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2119_wire : std_logic_vector(31 downto 0);
    signal type_cast_2122_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2128_wire : std_logic_vector(63 downto 0);
    signal type_cast_2145_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2150_wire : std_logic_vector(31 downto 0);
    signal type_cast_2153_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2159_wire : std_logic_vector(63 downto 0);
    signal type_cast_2175_wire : std_logic_vector(31 downto 0);
    signal type_cast_2181_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2199_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2207_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2212_wire : std_logic_vector(31 downto 0);
    signal type_cast_2230_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2236_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2248_wire : std_logic_vector(15 downto 0);
    signal type_cast_2250_wire : std_logic_vector(15 downto 0);
    signal type_cast_2254_wire : std_logic_vector(15 downto 0);
    signal type_cast_2256_wire : std_logic_vector(15 downto 0);
    signal type_cast_2260_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1879_word_address_0 <= "0";
    array_obj_ref_2135_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2135_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2135_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2135_resized_base_address <= "00000000000000";
    array_obj_ref_2166_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2166_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2166_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2166_resized_base_address <= "00000000000000";
    iNsTr_10_1942 <= "00000000000000000000000000000010";
    iNsTr_2_1825 <= "00000000000000000000000000000011";
    iNsTr_3_1847 <= "00000000000000000000000000000100";
    iNsTr_4_1857 <= "00000000000000000000000000000000";
    iNsTr_5_1873 <= "00000000000000000000000000000011";
    iNsTr_6_1890 <= "00000000000000000000000000000001";
    iNsTr_7_1906 <= "00000000000000000000000000000100";
    iNsTr_8_1918 <= "00000000000000000000000000000100";
    iNsTr_9_1930 <= "00000000000000000000000000000011";
    ptr_deref_1828_word_offset_0 <= "0000000";
    ptr_deref_1850_word_offset_0 <= "0000000";
    ptr_deref_1860_word_offset_0 <= "0";
    ptr_deref_1876_word_offset_0 <= "0000000";
    ptr_deref_1893_word_offset_0 <= "0";
    ptr_deref_1909_word_offset_0 <= "0000000";
    ptr_deref_1921_word_offset_0 <= "0000000";
    ptr_deref_1933_word_offset_0 <= "0000000";
    ptr_deref_1945_word_offset_0 <= "0000000";
    ptr_deref_2140_word_offset_0 <= "00000000000000";
    ptr_deref_2170_word_offset_0 <= "00000000000000";
    type_cast_1833_wire_constant <= "00000000000000000000000000000001";
    type_cast_1950_wire_constant <= "00000000000000000000000000000001";
    type_cast_1967_wire_constant <= "0000000000000000";
    type_cast_2027_wire_constant <= "00000000000000000000000000010000";
    type_cast_2033_wire_constant <= "11111111111111110000000000000000";
    type_cast_2041_wire_constant <= "00000000000000000000000000010000";
    type_cast_2048_wire_constant <= "00000000000000000000000000010000";
    type_cast_2054_wire_constant <= "11111111111111110000000000000000";
    type_cast_2062_wire_constant <= "00000000000000000000000000010000";
    type_cast_2089_wire_constant <= "0000000000000000";
    type_cast_2094_wire_constant <= "0000000000000100";
    type_cast_2114_wire_constant <= "00000000000000000000000000010000";
    type_cast_2122_wire_constant <= "00000000000000000000000000010010";
    type_cast_2145_wire_constant <= "00000000000000000000000000010000";
    type_cast_2153_wire_constant <= "00000000000000000000000000010010";
    type_cast_2181_wire_constant <= "00000000000000000000000000000100";
    type_cast_2199_wire_constant <= "0000000000000001";
    type_cast_2207_wire_constant <= "0000000000000001";
    type_cast_2230_wire_constant <= "0000000000000001";
    type_cast_2236_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1955: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1958_wire & type_cast_1960_wire;
      req <= phi_stmt_1955_req_0 & phi_stmt_1955_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1955",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1955_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1955,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1955
    phi_stmt_1961: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1964_wire & type_cast_1967_wire_constant;
      req <= phi_stmt_1961_req_0 & phi_stmt_1961_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1961",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1961_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1961,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1961
    phi_stmt_2083: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2086_wire & type_cast_2089_wire_constant;
      req <= phi_stmt_2083_req_0 & phi_stmt_2083_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2083",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2083_ack_0,
          idata => idata,
          odata => indvar_2083,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2083
    phi_stmt_2245: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2248_wire & type_cast_2250_wire;
      req <= phi_stmt_2245_req_0 & phi_stmt_2245_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2245",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2245_ack_0,
          idata => idata,
          odata => input_dim1x_x2_2245,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2245
    phi_stmt_2251: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2254_wire & type_cast_2256_wire;
      req <= phi_stmt_2251_req_0 & phi_stmt_2251_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2251",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2251_ack_0,
          idata => idata,
          odata => input_dim0x_x0_2251,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2251
    addr_of_2136_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2136_final_reg_req_0;
      addr_of_2136_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2136_final_reg_req_1;
      addr_of_2136_final_reg_ack_1<= rack(0);
      addr_of_2136_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2136_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2135_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2137,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2167_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2167_final_reg_req_0;
      addr_of_2167_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2167_final_reg_req_1;
      addr_of_2167_final_reg_ack_1<= rack(0);
      addr_of_2167_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2167_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2166_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx62_2168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1838_inst_req_0;
      type_cast_1838_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1838_inst_req_1;
      type_cast_1838_inst_ack_1<= rack(0);
      type_cast_1838_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1835,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1839,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1864_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1864_inst_req_0;
      type_cast_1864_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1864_inst_req_1;
      type_cast_1864_inst_ack_1<= rack(0);
      type_cast_1864_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1864_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp21_1861,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1865,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1883_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1883_inst_req_0;
      type_cast_1883_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1883_inst_req_1;
      type_cast_1883_inst_ack_1<= rack(0);
      type_cast_1883_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1883_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26_1880,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_1884,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1897_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1897_inst_req_0;
      type_cast_1897_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1897_inst_req_1;
      type_cast_1897_inst_ack_1<= rack(0);
      type_cast_1897_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1897_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp32_1894,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_1898,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1958_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1958_inst_req_0;
      type_cast_1958_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1958_inst_req_1;
      type_cast_1958_inst_ack_1<= rack(0);
      type_cast_1958_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1958_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_1839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1958_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1960_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1960_inst_req_0;
      type_cast_1960_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1960_inst_req_1;
      type_cast_1960_inst_ack_1<= rack(0);
      type_cast_1960_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1960_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1960_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1964_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1964_inst_req_0;
      type_cast_1964_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1964_inst_req_1;
      type_cast_1964_inst_ack_1<= rack(0);
      type_cast_1964_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1964_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1964_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1972_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1972_inst_req_0;
      type_cast_1972_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1972_inst_req_1;
      type_cast_1972_inst_ack_1<= rack(0);
      type_cast_1972_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1972_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1971_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1973,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1977_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1977_inst_req_0;
      type_cast_1977_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1977_inst_req_1;
      type_cast_1977_inst_ack_1<= rack(0);
      type_cast_1977_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1977_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1976_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_1978,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2038_inst
    process(sext_2035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2035(31 downto 0);
      type_cast_2038_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2043_inst
    process(ASHR_i32_i32_2042_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2042_wire(31 downto 0);
      conv46_2044 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2059_inst
    process(sext103_2056) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext103_2056(31 downto 0);
      type_cast_2059_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2064_inst
    process(ASHR_i32_i32_2063_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2063_wire(31 downto 0);
      conv49_2065 <= tmp_var; -- 
    end process;
    type_cast_2086_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2086_inst_req_0;
      type_cast_2086_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2086_inst_req_1;
      type_cast_2086_inst_ack_1<= rack(0);
      type_cast_2086_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2086_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2201,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2086_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2099_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2099_inst_req_0;
      type_cast_2099_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2099_inst_req_1;
      type_cast_2099_inst_ack_1<= rack(0);
      type_cast_2099_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2099_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2096,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9102_2100,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2119_inst
    process(sext105_2116) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext105_2116(31 downto 0);
      type_cast_2119_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2124_inst
    process(ASHR_i32_i32_2123_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2123_wire(31 downto 0);
      shr_2125 <= tmp_var; -- 
    end process;
    type_cast_2129_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2129_inst_req_0;
      type_cast_2129_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2129_inst_req_1;
      type_cast_2129_inst_ack_1<= rack(0);
      type_cast_2129_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2129_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2128_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2130,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2150_inst
    process(sext106_2147) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext106_2147(31 downto 0);
      type_cast_2150_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2155_inst
    process(ASHR_i32_i32_2154_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2154_wire(31 downto 0);
      shr60_2156 <= tmp_var; -- 
    end process;
    type_cast_2160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2160_inst_req_0;
      type_cast_2160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2160_inst_req_1;
      type_cast_2160_inst_ack_1<= rack(0);
      type_cast_2160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2159_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom61_2161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2176_inst_req_0;
      type_cast_2176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2176_inst_req_1;
      type_cast_2176_inst_ack_1<= rack(0);
      type_cast_2176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2175_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2213_inst_req_0;
      type_cast_2213_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2213_inst_req_1;
      type_cast_2213_inst_ack_1<= rack(0);
      type_cast_2213_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2213_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2212_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2214,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2241_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2241_inst_req_0;
      type_cast_2241_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2241_inst_req_1;
      type_cast_2241_inst_ack_1<= rack(0);
      type_cast_2241_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2241_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div83_2238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_2242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2248_inst_req_0;
      type_cast_2248_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2248_inst_req_1;
      type_cast_2248_inst_ack_1<= rack(0);
      type_cast_2248_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2248_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_2209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2248_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2250_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2250_inst_req_0;
      type_cast_2250_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2250_inst_req_1;
      type_cast_2250_inst_ack_1<= rack(0);
      type_cast_2250_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2250_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv84_2242,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2250_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2254_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2254_inst_req_0;
      type_cast_2254_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2254_inst_req_1;
      type_cast_2254_inst_ack_1<= rack(0);
      type_cast_2254_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2254_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc81_2232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2254_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2256_inst_req_0;
      type_cast_2256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2256_inst_req_1;
      type_cast_2256_inst_ack_1<= rack(0);
      type_cast_2256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2x_xph_1961,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2256_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2261_inst_req_0;
      type_cast_2261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2261_inst_req_1;
      type_cast_2261_inst_ack_1<= rack(0);
      type_cast_2261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2260_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_2262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1879_gather_scatter
    process(LOAD_padding_1879_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1879_data_0;
      ov(15 downto 0) := iv;
      tmp26_1880 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2135_index_1_rename
    process(R_idxprom_2134_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2134_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2134_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2135_index_1_resize
    process(idxprom_2130) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2130;
      ov := iv(13 downto 0);
      R_idxprom_2134_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2135_root_address_inst
    process(array_obj_ref_2135_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2135_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2135_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2166_index_1_rename
    process(R_idxprom61_2165_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom61_2165_resized;
      ov(13 downto 0) := iv;
      R_idxprom61_2165_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2166_index_1_resize
    process(idxprom61_2161) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom61_2161;
      ov := iv(13 downto 0);
      R_idxprom61_2165_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2166_root_address_inst
    process(array_obj_ref_2166_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2166_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2166_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1828_addr_0
    process(ptr_deref_1828_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1828_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1828_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1828_base_resize
    process(iNsTr_2_1825) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1825;
      ov := iv(6 downto 0);
      ptr_deref_1828_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1828_gather_scatter
    process(ptr_deref_1828_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1828_data_0;
      ov(31 downto 0) := iv;
      tmp_1829 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1828_root_address_inst
    process(ptr_deref_1828_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1828_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1828_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1850_addr_0
    process(ptr_deref_1850_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1850_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1850_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1850_base_resize
    process(iNsTr_3_1847) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1847;
      ov := iv(6 downto 0);
      ptr_deref_1850_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1850_gather_scatter
    process(ptr_deref_1850_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1850_data_0;
      ov(31 downto 0) := iv;
      tmp10_1851 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1850_root_address_inst
    process(ptr_deref_1850_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1850_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1850_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1860_addr_0
    process(ptr_deref_1860_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1860_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1860_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1860_base_resize
    process(iNsTr_4_1857) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1857;
      ov := iv(0 downto 0);
      ptr_deref_1860_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1860_gather_scatter
    process(ptr_deref_1860_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1860_data_0;
      ov(15 downto 0) := iv;
      tmp21_1861 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1860_root_address_inst
    process(ptr_deref_1860_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1860_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1860_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1876_addr_0
    process(ptr_deref_1876_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1876_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1876_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1876_base_resize
    process(iNsTr_5_1873) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1873;
      ov := iv(6 downto 0);
      ptr_deref_1876_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1876_gather_scatter
    process(ptr_deref_1876_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1876_data_0;
      ov(31 downto 0) := iv;
      tmp24_1877 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1876_root_address_inst
    process(ptr_deref_1876_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1876_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1876_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1893_addr_0
    process(ptr_deref_1893_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1893_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1893_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1893_base_resize
    process(iNsTr_6_1890) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1890;
      ov := iv(0 downto 0);
      ptr_deref_1893_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1893_gather_scatter
    process(ptr_deref_1893_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1893_data_0;
      ov(15 downto 0) := iv;
      tmp32_1894 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1893_root_address_inst
    process(ptr_deref_1893_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1893_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1893_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1909_addr_0
    process(ptr_deref_1909_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1909_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1909_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1909_base_resize
    process(iNsTr_7_1906) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1906;
      ov := iv(6 downto 0);
      ptr_deref_1909_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1909_gather_scatter
    process(ptr_deref_1909_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1909_data_0;
      ov(31 downto 0) := iv;
      tmp35_1910 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1909_root_address_inst
    process(ptr_deref_1909_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1909_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1909_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1921_addr_0
    process(ptr_deref_1921_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1921_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1921_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1921_base_resize
    process(iNsTr_8_1918) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1918;
      ov := iv(6 downto 0);
      ptr_deref_1921_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1921_gather_scatter
    process(ptr_deref_1921_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1921_data_0;
      ov(31 downto 0) := iv;
      tmp44_1922 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1921_root_address_inst
    process(ptr_deref_1921_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1921_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1921_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1933_addr_0
    process(ptr_deref_1933_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1933_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1933_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1933_base_resize
    process(iNsTr_9_1930) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1930;
      ov := iv(6 downto 0);
      ptr_deref_1933_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1933_gather_scatter
    process(ptr_deref_1933_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1933_data_0;
      ov(31 downto 0) := iv;
      tmp47_1934 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1933_root_address_inst
    process(ptr_deref_1933_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1933_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1933_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1945_addr_0
    process(ptr_deref_1945_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1945_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1945_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1945_base_resize
    process(iNsTr_10_1942) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1942;
      ov := iv(6 downto 0);
      ptr_deref_1945_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1945_gather_scatter
    process(ptr_deref_1945_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1945_data_0;
      ov(31 downto 0) := iv;
      tmp87_1946 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1945_root_address_inst
    process(ptr_deref_1945_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1945_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1945_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2140_addr_0
    process(ptr_deref_2140_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2140_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2140_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2140_base_resize
    process(arrayidx_2137) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2137;
      ov := iv(13 downto 0);
      ptr_deref_2140_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2140_gather_scatter
    process(ptr_deref_2140_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2140_data_0;
      ov(63 downto 0) := iv;
      tmp57_2141 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2140_root_address_inst
    process(ptr_deref_2140_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2140_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2140_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2170_addr_0
    process(ptr_deref_2170_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2170_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2170_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2170_base_resize
    process(arrayidx62_2168) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx62_2168;
      ov := iv(13 downto 0);
      ptr_deref_2170_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2170_gather_scatter
    process(tmp57_2141) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp57_2141;
      ov(63 downto 0) := iv;
      ptr_deref_2170_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2170_root_address_inst
    process(ptr_deref_2170_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2170_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2170_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2189_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2188;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2189_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2189_branch_req_0,
          ack0 => if_stmt_2189_branch_ack_0,
          ack1 => if_stmt_2189_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2220_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_2219;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2220_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2220_branch_req_0,
          ack0 => if_stmt_2220_branch_ack_0,
          ack1 => if_stmt_2220_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2268_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp89_2267;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2268_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2268_branch_req_0,
          ack0 => if_stmt_2268_branch_ack_0,
          ack1 => if_stmt_2268_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2200_inst
    process(indvar_2083) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2083, type_cast_2199_wire_constant, tmp_var);
      indvarx_xnext_2201 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2208_inst
    process(input_dim1x_x1x_xph_1955) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1955, type_cast_2207_wire_constant, tmp_var);
      inc_2209 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2231_inst
    process(input_dim0x_x2x_xph_1961) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_1961, type_cast_2230_wire_constant, tmp_var);
      inc81_2232 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1987_inst
    process(mul_1983, conv12_1973) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_1983, conv12_1973, tmp_var);
      add_1988 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2002_inst
    process(mul23_1998, tmp24_1877) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul23_1998, tmp24_1877, tmp_var);
      add25_2003 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2017_inst
    process(mul34_2013, tmp35_1910) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul34_2013, tmp35_1910, tmp_var);
      add36_2018 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2034_inst
    process(sub40_2029) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub40_2029, type_cast_2033_wire_constant, tmp_var);
      sext_2035 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2055_inst
    process(sub28_2050) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub28_2050, type_cast_2054_wire_constant, tmp_var);
      sext103_2056 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2074_inst
    process(conv46_2044, mul50_2070) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv46_2044, mul50_2070, tmp_var);
      add51_2075 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2104_inst
    process(mul16_1993, conv9102_2100) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul16_1993, conv9102_2100, tmp_var);
      add17_2105 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2109_inst
    process(mul52_2080, conv9102_2100) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul52_2080, conv9102_2100, tmp_var);
      add53_2110 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2182_inst
    process(conv65_2177) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv65_2177, type_cast_2181_wire_constant, tmp_var);
      add66_2183 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2042_inst
    process(type_cast_2038_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2038_wire, type_cast_2041_wire_constant, tmp_var);
      ASHR_i32_i32_2042_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2063_inst
    process(type_cast_2059_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2059_wire, type_cast_2062_wire_constant, tmp_var);
      ASHR_i32_i32_2063_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2123_inst
    process(type_cast_2119_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2119_wire, type_cast_2122_wire_constant, tmp_var);
      ASHR_i32_i32_2123_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2154_inst
    process(type_cast_2150_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2150_wire, type_cast_2153_wire_constant, tmp_var);
      ASHR_i32_i32_2154_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2218_inst
    process(conv75_2214, tmp_1829) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv75_2214, tmp_1829, tmp_var);
      cmp77_2219 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2266_inst
    process(conv86_2262, div88_1952) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv86_2262, div88_1952, tmp_var);
      cmp89_2267 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1834_inst
    process(tmp_1829) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1829, type_cast_1833_wire_constant, tmp_var);
      div_1835 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1951_inst
    process(tmp87_1946) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp87_1946, type_cast_1950_wire_constant, tmp_var);
      div88_1952 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2237_inst
    process(tmp_1829) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1829, type_cast_2236_wire_constant, tmp_var);
      div83_2238 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2095_inst
    process(indvar_2083) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2083, type_cast_2094_wire_constant, tmp_var);
      input_dim2x_x1_2096 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1982_inst
    process(tmp_1829, conv15_1978) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1829, conv15_1978, tmp_var);
      mul_1983 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1992_inst
    process(add_1988, tmp10_1851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1988, tmp10_1851, tmp_var);
      mul16_1993 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1997_inst
    process(conv22_1865, conv15_1978) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv22_1865, conv15_1978, tmp_var);
      mul23_1998 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2012_inst
    process(conv33_1898, conv12_1973) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv33_1898, conv12_1973, tmp_var);
      mul34_2013 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2069_inst
    process(tmp47_1934, conv49_2065) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp47_1934, conv49_2065, tmp_var);
      mul50_2070 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2079_inst
    process(add51_2075, tmp44_1922) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add51_2075, tmp44_1922, tmp_var);
      mul52_2080 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2028_inst
    process(sub39_2023) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub39_2023, type_cast_2027_wire_constant, tmp_var);
      sub40_2029 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2049_inst
    process(sub_2008) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2008, type_cast_2048_wire_constant, tmp_var);
      sub28_2050 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2115_inst
    process(add17_2105) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add17_2105, type_cast_2114_wire_constant, tmp_var);
      sext105_2116 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2146_inst
    process(add53_2110) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add53_2110, type_cast_2145_wire_constant, tmp_var);
      sext106_2147 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2007_inst
    process(add25_2003, conv27_1884) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add25_2003, conv27_1884, tmp_var);
      sub_2008 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2022_inst
    process(add36_2018, conv27_1884) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add36_2018, conv27_1884, tmp_var);
      sub39_2023 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2187_inst
    process(add66_2183, tmp10_1851) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add66_2183, tmp10_1851, tmp_var);
      cmp_2188 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_2135_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2134_scaled;
      array_obj_ref_2135_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2135_index_offset_req_0;
      array_obj_ref_2135_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2135_index_offset_req_1;
      array_obj_ref_2135_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_2166_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom61_2165_scaled;
      array_obj_ref_2166_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2166_index_offset_req_0;
      array_obj_ref_2166_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2166_index_offset_req_1;
      array_obj_ref_2166_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- unary operator type_cast_1971_inst
    process(input_dim1x_x1x_xph_1955) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_1955, tmp_var);
      type_cast_1971_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1976_inst
    process(input_dim0x_x2x_xph_1961) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_1961, tmp_var);
      type_cast_1976_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2128_inst
    process(shr_2125) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2125, tmp_var);
      type_cast_2128_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2159_inst
    process(shr60_2156) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr60_2156, tmp_var);
      type_cast_2159_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2175_inst
    process(input_dim2x_x1_2096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2096, tmp_var);
      type_cast_2175_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2212_inst
    process(inc_2209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2209, tmp_var);
      type_cast_2212_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2260_inst
    process(input_dim0x_x0_2251) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_2251, tmp_var);
      type_cast_2260_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1879_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1879_load_0_req_0;
      LOAD_padding_1879_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1879_load_0_req_1;
      LOAD_padding_1879_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1879_word_address_0;
      LOAD_padding_1879_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1945_load_0 ptr_deref_1850_load_0 ptr_deref_1828_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1945_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1850_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1828_load_0_req_0;
      ptr_deref_1945_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1850_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1828_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1945_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1850_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1828_load_0_req_1;
      ptr_deref_1945_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1850_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1828_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1945_word_address_0 & ptr_deref_1850_word_address_0 & ptr_deref_1828_word_address_0;
      ptr_deref_1945_data_0 <= data_out(95 downto 64);
      ptr_deref_1850_data_0 <= data_out(63 downto 32);
      ptr_deref_1828_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1893_load_0 ptr_deref_1860_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1893_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1860_load_0_req_0;
      ptr_deref_1893_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1860_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1893_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1860_load_0_req_1;
      ptr_deref_1893_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1860_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1893_word_address_0 & ptr_deref_1860_word_address_0;
      ptr_deref_1893_data_0 <= data_out(31 downto 16);
      ptr_deref_1860_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1876_load_0 ptr_deref_1909_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1876_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1909_load_0_req_0;
      ptr_deref_1876_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1909_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1876_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1909_load_0_req_1;
      ptr_deref_1876_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1909_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1876_word_address_0 & ptr_deref_1909_word_address_0;
      ptr_deref_1876_data_0 <= data_out(63 downto 32);
      ptr_deref_1909_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1921_load_0 ptr_deref_1933_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1921_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1933_load_0_req_0;
      ptr_deref_1921_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1933_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1921_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1933_load_0_req_1;
      ptr_deref_1921_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1933_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1921_word_address_0 & ptr_deref_1933_word_address_0;
      ptr_deref_1921_data_0 <= data_out(63 downto 32);
      ptr_deref_1933_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2140_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2140_load_0_req_0;
      ptr_deref_2140_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2140_load_0_req_1;
      ptr_deref_2140_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2140_word_address_0;
      ptr_deref_2140_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2170_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2170_store_0_req_0;
      ptr_deref_2170_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2170_store_0_req_1;
      ptr_deref_2170_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2170_word_address_0;
      data_in <= ptr_deref_2170_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1815_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_start_1815_inst_req_0;
      RPIPE_Block1_start_1815_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_start_1815_inst_req_1;
      RPIPE_Block1_start_1815_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1816 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2276_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2276_inst_req_0;
      WPIPE_Block1_done_2276_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2276_inst_req_1;
      WPIPE_Block1_done_2276_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1816;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_6511_start: Boolean;
  signal convTransposeC_CP_6511_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_2299_load_0_ack_1 : boolean;
  signal type_cast_2647_inst_req_1 : boolean;
  signal type_cast_2647_inst_ack_0 : boolean;
  signal type_cast_2438_inst_req_0 : boolean;
  signal ptr_deref_2299_load_0_req_0 : boolean;
  signal ptr_deref_2299_load_0_ack_0 : boolean;
  signal type_cast_2309_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2286_inst_req_1 : boolean;
  signal phi_stmt_2433_req_1 : boolean;
  signal type_cast_2309_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2286_inst_ack_1 : boolean;
  signal type_cast_2647_inst_req_0 : boolean;
  signal type_cast_2309_inst_ack_1 : boolean;
  signal type_cast_2560_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2286_inst_req_0 : boolean;
  signal ptr_deref_2299_load_0_req_1 : boolean;
  signal type_cast_2647_inst_ack_1 : boolean;
  signal if_stmt_2660_branch_ack_0 : boolean;
  signal type_cast_2438_inst_ack_1 : boolean;
  signal ptr_deref_2321_load_0_req_0 : boolean;
  signal ptr_deref_2321_load_0_req_1 : boolean;
  signal WPIPE_Block2_done_2725_inst_ack_1 : boolean;
  signal ptr_deref_2321_load_0_ack_1 : boolean;
  signal WPIPE_Block2_done_2725_inst_req_1 : boolean;
  signal type_cast_2560_inst_req_0 : boolean;
  signal ptr_deref_2321_load_0_ack_0 : boolean;
  signal RPIPE_Block2_start_2286_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2725_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2725_inst_req_0 : boolean;
  signal ptr_deref_2641_store_0_ack_1 : boolean;
  signal ptr_deref_2641_store_0_req_1 : boolean;
  signal type_cast_2309_inst_ack_0 : boolean;
  signal ptr_deref_2333_load_0_req_0 : boolean;
  signal ptr_deref_2333_load_0_ack_0 : boolean;
  signal type_cast_2432_inst_req_0 : boolean;
  signal ptr_deref_2641_store_0_ack_0 : boolean;
  signal addr_of_2638_final_reg_req_1 : boolean;
  signal if_stmt_2660_branch_ack_1 : boolean;
  signal if_stmt_2717_branch_ack_0 : boolean;
  signal if_stmt_2717_branch_ack_1 : boolean;
  signal if_stmt_2717_branch_req_0 : boolean;
  signal ptr_deref_2333_load_0_req_1 : boolean;
  signal ptr_deref_2333_load_0_ack_1 : boolean;
  signal addr_of_2638_final_reg_ack_1 : boolean;
  signal type_cast_2438_inst_req_1 : boolean;
  signal type_cast_2432_inst_ack_0 : boolean;
  signal phi_stmt_2426_req_0 : boolean;
  signal phi_stmt_2426_ack_0 : boolean;
  signal ptr_deref_2343_load_0_req_0 : boolean;
  signal ptr_deref_2343_load_0_ack_0 : boolean;
  signal ptr_deref_2343_load_0_req_1 : boolean;
  signal type_cast_2710_inst_ack_1 : boolean;
  signal ptr_deref_2343_load_0_ack_1 : boolean;
  signal type_cast_2710_inst_req_1 : boolean;
  signal phi_stmt_2433_req_0 : boolean;
  signal ptr_deref_2641_store_0_req_0 : boolean;
  signal phi_stmt_2426_req_1 : boolean;
  signal type_cast_2710_inst_ack_0 : boolean;
  signal type_cast_2436_inst_ack_1 : boolean;
  signal type_cast_2347_inst_req_0 : boolean;
  signal type_cast_2436_inst_req_1 : boolean;
  signal type_cast_2347_inst_ack_0 : boolean;
  signal addr_of_2638_final_reg_ack_0 : boolean;
  signal type_cast_2347_inst_req_1 : boolean;
  signal type_cast_2347_inst_ack_1 : boolean;
  signal type_cast_2432_inst_ack_1 : boolean;
  signal type_cast_2432_inst_req_1 : boolean;
  signal type_cast_2436_inst_ack_0 : boolean;
  signal type_cast_2436_inst_req_0 : boolean;
  signal ptr_deref_2359_load_0_req_0 : boolean;
  signal ptr_deref_2359_load_0_ack_0 : boolean;
  signal if_stmt_2660_branch_req_0 : boolean;
  signal ptr_deref_2359_load_0_req_1 : boolean;
  signal type_cast_2710_inst_req_0 : boolean;
  signal ptr_deref_2359_load_0_ack_1 : boolean;
  signal addr_of_2638_final_reg_req_0 : boolean;
  signal type_cast_2693_inst_ack_1 : boolean;
  signal LOAD_padding_2362_load_0_req_0 : boolean;
  signal type_cast_2693_inst_req_1 : boolean;
  signal LOAD_padding_2362_load_0_ack_0 : boolean;
  signal LOAD_padding_2362_load_0_req_1 : boolean;
  signal LOAD_padding_2362_load_0_ack_1 : boolean;
  signal type_cast_2693_inst_ack_0 : boolean;
  signal type_cast_2438_inst_ack_0 : boolean;
  signal type_cast_2693_inst_req_0 : boolean;
  signal type_cast_2366_inst_req_0 : boolean;
  signal type_cast_2366_inst_ack_0 : boolean;
  signal type_cast_2366_inst_req_1 : boolean;
  signal type_cast_2366_inst_ack_1 : boolean;
  signal type_cast_2684_inst_ack_1 : boolean;
  signal type_cast_2684_inst_req_1 : boolean;
  signal type_cast_2684_inst_ack_0 : boolean;
  signal type_cast_2684_inst_req_0 : boolean;
  signal ptr_deref_2376_load_0_req_0 : boolean;
  signal ptr_deref_2376_load_0_ack_0 : boolean;
  signal ptr_deref_2376_load_0_req_1 : boolean;
  signal ptr_deref_2376_load_0_ack_1 : boolean;
  signal type_cast_2380_inst_req_0 : boolean;
  signal type_cast_2380_inst_ack_0 : boolean;
  signal type_cast_2380_inst_req_1 : boolean;
  signal type_cast_2380_inst_ack_1 : boolean;
  signal ptr_deref_2392_load_0_req_0 : boolean;
  signal ptr_deref_2392_load_0_ack_0 : boolean;
  signal ptr_deref_2392_load_0_req_1 : boolean;
  signal ptr_deref_2392_load_0_ack_1 : boolean;
  signal ptr_deref_2404_load_0_req_0 : boolean;
  signal ptr_deref_2404_load_0_ack_0 : boolean;
  signal ptr_deref_2404_load_0_req_1 : boolean;
  signal ptr_deref_2404_load_0_ack_1 : boolean;
  signal ptr_deref_2416_load_0_req_0 : boolean;
  signal ptr_deref_2416_load_0_ack_0 : boolean;
  signal ptr_deref_2416_load_0_req_1 : boolean;
  signal ptr_deref_2416_load_0_ack_1 : boolean;
  signal type_cast_2443_inst_req_0 : boolean;
  signal type_cast_2443_inst_ack_0 : boolean;
  signal type_cast_2443_inst_req_1 : boolean;
  signal type_cast_2443_inst_ack_1 : boolean;
  signal type_cast_2448_inst_req_0 : boolean;
  signal type_cast_2448_inst_ack_0 : boolean;
  signal type_cast_2448_inst_req_1 : boolean;
  signal type_cast_2448_inst_ack_1 : boolean;
  signal type_cast_2570_inst_req_0 : boolean;
  signal type_cast_2570_inst_ack_0 : boolean;
  signal type_cast_2570_inst_req_1 : boolean;
  signal type_cast_2570_inst_ack_1 : boolean;
  signal type_cast_2600_inst_req_0 : boolean;
  signal type_cast_2600_inst_ack_0 : boolean;
  signal type_cast_2600_inst_req_1 : boolean;
  signal type_cast_2600_inst_ack_1 : boolean;
  signal array_obj_ref_2606_index_offset_req_0 : boolean;
  signal array_obj_ref_2606_index_offset_ack_0 : boolean;
  signal array_obj_ref_2606_index_offset_req_1 : boolean;
  signal array_obj_ref_2606_index_offset_ack_1 : boolean;
  signal addr_of_2607_final_reg_req_0 : boolean;
  signal addr_of_2607_final_reg_ack_0 : boolean;
  signal addr_of_2607_final_reg_req_1 : boolean;
  signal addr_of_2607_final_reg_ack_1 : boolean;
  signal phi_stmt_2433_ack_0 : boolean;
  signal ptr_deref_2611_load_0_req_0 : boolean;
  signal ptr_deref_2611_load_0_ack_0 : boolean;
  signal ptr_deref_2611_load_0_req_1 : boolean;
  signal ptr_deref_2611_load_0_ack_1 : boolean;
  signal type_cast_2631_inst_req_0 : boolean;
  signal type_cast_2631_inst_ack_0 : boolean;
  signal type_cast_2631_inst_req_1 : boolean;
  signal type_cast_2631_inst_ack_1 : boolean;
  signal array_obj_ref_2637_index_offset_req_0 : boolean;
  signal array_obj_ref_2637_index_offset_ack_0 : boolean;
  signal array_obj_ref_2637_index_offset_req_1 : boolean;
  signal array_obj_ref_2637_index_offset_ack_1 : boolean;
  signal type_cast_2560_inst_req_1 : boolean;
  signal type_cast_2560_inst_ack_1 : boolean;
  signal phi_stmt_2554_req_1 : boolean;
  signal phi_stmt_2554_req_0 : boolean;
  signal phi_stmt_2554_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_6511_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6511_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_6511_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6511_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_6511: Block -- control-path 
    signal convTransposeC_CP_6511_elements: BooleanArray(92 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_6511_elements(0) <= convTransposeC_CP_6511_start;
    convTransposeC_CP_6511_symbol <= convTransposeC_CP_6511_elements(70);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2284/assign_stmt_2287/$entry
      -- CP-element group 0: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2284/assign_stmt_2287__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2284/branch_block_stmt_2284__entry__
      -- CP-element group 0: 	 branch_block_stmt_2284/$entry
      -- CP-element group 0: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_Sample/$entry
      -- 
    rr_6559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(0), ack => RPIPE_Block2_start_2286_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_Sample/ra
      -- 
    ra_6560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2286_inst_ack_0, ack => convTransposeC_CP_6511_elements(1)); -- 
    cr_6564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(1), ack => RPIPE_Block2_start_2286_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2:  members (265) 
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2287/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2287__exit__
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2287/RPIPE_Block2_start_2286_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423__entry__
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/word_access_complete/word_0/cr
      -- 
    ca_6565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2286_inst_ack_1, ack => convTransposeC_CP_6511_elements(2)); -- 
    rr_6601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2299_load_0_req_0); -- 
    cr_6631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => type_cast_2309_inst_req_1); -- 
    cr_6612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2299_load_0_req_1); -- 
    rr_6665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2321_load_0_req_0); -- 
    cr_6676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2321_load_0_req_1); -- 
    rr_6715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2333_load_0_req_0); -- 
    cr_6726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2333_load_0_req_1); -- 
    rr_6765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2343_load_0_req_0); -- 
    cr_6776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2343_load_0_req_1); -- 
    cr_6795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => type_cast_2347_inst_req_1); -- 
    rr_6829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2359_load_0_req_0); -- 
    cr_6840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2359_load_0_req_1); -- 
    rr_6862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => LOAD_padding_2362_load_0_req_0); -- 
    cr_6873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => LOAD_padding_2362_load_0_req_1); -- 
    cr_6892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => type_cast_2366_inst_req_1); -- 
    rr_6926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2376_load_0_req_0); -- 
    cr_6937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2376_load_0_req_1); -- 
    cr_6956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => type_cast_2380_inst_req_1); -- 
    rr_6990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2392_load_0_req_0); -- 
    cr_7001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2392_load_0_req_1); -- 
    rr_7040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2404_load_0_req_0); -- 
    cr_7051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2404_load_0_req_1); -- 
    rr_7090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2416_load_0_req_0); -- 
    cr_7101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2416_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_sample_completed_
      -- 
    ra_6602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2299_load_0_ack_0, ack => convTransposeC_CP_6511_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/ptr_deref_2299_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/ptr_deref_2299_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/ptr_deref_2299_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2299_Update/ptr_deref_2299_Merge/$entry
      -- 
    ca_6613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2299_load_0_ack_1, ack => convTransposeC_CP_6511_elements(4)); -- 
    rr_6626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(4), ack => type_cast_2309_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_Sample/ra
      -- 
    ra_6627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_0, ack => convTransposeC_CP_6511_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2309_update_completed_
      -- 
    ca_6632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_1, ack => convTransposeC_CP_6511_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_sample_completed_
      -- 
    ra_6666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2321_load_0_ack_0, ack => convTransposeC_CP_6511_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	31 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/ptr_deref_2321_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/ptr_deref_2321_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/ptr_deref_2321_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/ptr_deref_2321_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2321_Update/word_access_complete/word_0/$exit
      -- 
    ca_6677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2321_load_0_ack_1, ack => convTransposeC_CP_6511_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Sample/word_access_start/word_0/ra
      -- 
    ra_6716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2333_load_0_ack_0, ack => convTransposeC_CP_6511_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	31 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/ptr_deref_2333_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/ptr_deref_2333_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/ptr_deref_2333_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2333_Update/ptr_deref_2333_Merge/merge_ack
      -- 
    ca_6727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2333_load_0_ack_1, ack => convTransposeC_CP_6511_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Sample/word_access_start/word_0/ra
      -- 
    ra_6766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2343_load_0_ack_0, ack => convTransposeC_CP_6511_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (12) 
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/ptr_deref_2343_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/ptr_deref_2343_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/ptr_deref_2343_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2343_Update/ptr_deref_2343_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_Sample/rr
      -- 
    ca_6777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2343_load_0_ack_1, ack => convTransposeC_CP_6511_elements(12)); -- 
    rr_6790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(12), ack => type_cast_2347_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_Sample/ra
      -- 
    ra_6791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_0, ack => convTransposeC_CP_6511_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2347_Update/ca
      -- 
    ca_6796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_1, ack => convTransposeC_CP_6511_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Sample/word_access_start/word_0/ra
      -- 
    ra_6830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2359_load_0_ack_0, ack => convTransposeC_CP_6511_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/ptr_deref_2359_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/ptr_deref_2359_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/ptr_deref_2359_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2359_Update/ptr_deref_2359_Merge/merge_ack
      -- 
    ca_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2359_load_0_ack_1, ack => convTransposeC_CP_6511_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Sample/word_access_start/word_0/ra
      -- 
    ra_6863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2362_load_0_ack_0, ack => convTransposeC_CP_6511_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (12) 
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/LOAD_padding_2362_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/LOAD_padding_2362_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/LOAD_padding_2362_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/LOAD_padding_2362_Update/LOAD_padding_2362_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_Sample/rr
      -- 
    ca_6874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2362_load_0_ack_1, ack => convTransposeC_CP_6511_elements(18)); -- 
    rr_6887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(18), ack => type_cast_2366_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_Sample/ra
      -- 
    ra_6888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2366_inst_ack_0, ack => convTransposeC_CP_6511_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	31 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2366_Update/ca
      -- 
    ca_6893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2366_inst_ack_1, ack => convTransposeC_CP_6511_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Sample/word_access_start/word_0/ra
      -- 
    ra_6927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2376_load_0_ack_0, ack => convTransposeC_CP_6511_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (12) 
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/ptr_deref_2376_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/ptr_deref_2376_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/ptr_deref_2376_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2376_Update/ptr_deref_2376_Merge/merge_ack
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_Sample/rr
      -- 
    ca_6938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2376_load_0_ack_1, ack => convTransposeC_CP_6511_elements(22)); -- 
    rr_6951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(22), ack => type_cast_2380_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_Sample/ra
      -- 
    ra_6952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2380_inst_ack_0, ack => convTransposeC_CP_6511_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	31 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/type_cast_2380_Update/ca
      -- 
    ca_6957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2380_inst_ack_1, ack => convTransposeC_CP_6511_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Sample/word_access_start/word_0/ra
      -- 
    ra_6991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2392_load_0_ack_0, ack => convTransposeC_CP_6511_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/ptr_deref_2392_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/ptr_deref_2392_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/ptr_deref_2392_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2392_Update/ptr_deref_2392_Merge/merge_ack
      -- 
    ca_7002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2392_load_0_ack_1, ack => convTransposeC_CP_6511_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Sample/word_access_start/word_0/ra
      -- 
    ra_7041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_load_0_ack_0, ack => convTransposeC_CP_6511_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/ptr_deref_2404_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/ptr_deref_2404_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/ptr_deref_2404_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2404_Update/ptr_deref_2404_Merge/merge_ack
      -- 
    ca_7052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_load_0_ack_1, ack => convTransposeC_CP_6511_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Sample/word_access_start/word_0/ra
      -- 
    ra_7091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2416_load_0_ack_0, ack => convTransposeC_CP_6511_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/ptr_deref_2416_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/ptr_deref_2416_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/ptr_deref_2416_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/ptr_deref_2416_Update/ptr_deref_2416_Merge/merge_ack
      -- 
    ca_7102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2416_load_0_ack_1, ack => convTransposeC_CP_6511_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	8 
    -- CP-element group 31: 	24 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	10 
    -- CP-element group 31: 	20 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	6 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	72 
    -- CP-element group 31: 	73 
    -- CP-element group 31: 	71 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423__exit__
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/$entry
      -- CP-element group 31: 	 branch_block_stmt_2284/assign_stmt_2296_to_assign_stmt_2423/$exit
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/$entry
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/$entry
      -- 
    cr_7524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(31), ack => type_cast_2436_inst_req_1); -- 
    rr_7519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(31), ack => type_cast_2436_inst_req_0); -- 
    convTransposeC_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(16) & convTransposeC_CP_6511_elements(28) & convTransposeC_CP_6511_elements(8) & convTransposeC_CP_6511_elements(24) & convTransposeC_CP_6511_elements(14) & convTransposeC_CP_6511_elements(10) & convTransposeC_CP_6511_elements(20) & convTransposeC_CP_6511_elements(26) & convTransposeC_CP_6511_elements(30) & convTransposeC_CP_6511_elements(6);
      gj_convTransposeC_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	86 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_Sample/ra
      -- 
    ra_7119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2443_inst_ack_0, ack => convTransposeC_CP_6511_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	86 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_Update/ca
      -- 
    ca_7124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2443_inst_ack_1, ack => convTransposeC_CP_6511_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	86 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_Sample/ra
      -- 
    ra_7133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2448_inst_ack_0, ack => convTransposeC_CP_6511_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	86 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_Update/ca
      -- 
    ca_7138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2448_inst_ack_1, ack => convTransposeC_CP_6511_elements(35)); -- 
    -- CP-element group 36:  join  transition  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: 	33 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	90 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_2284/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 36: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551__exit__
      -- CP-element group 36: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/$exit
      -- CP-element group 36: 	 branch_block_stmt_2284/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_2284/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2554/$entry
      -- CP-element group 36: 	 branch_block_stmt_2284/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/$entry
      -- 
    convTransposeC_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(35) & convTransposeC_CP_6511_elements(33);
      gj_convTransposeC_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_Sample/ra
      -- 
    ra_7150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2570_inst_ack_0, ack => convTransposeC_CP_6511_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	92 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	47 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_Sample/rr
      -- 
    ca_7155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2570_inst_ack_1, ack => convTransposeC_CP_6511_elements(38)); -- 
    rr_7163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(38), ack => type_cast_2600_inst_req_0); -- 
    rr_7273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(38), ack => type_cast_2631_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_Sample/ra
      -- 
    ra_7164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2600_inst_ack_0, ack => convTransposeC_CP_6511_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	92 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (16) 
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_resized_1
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_scaled_1
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_computed_1
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_resize_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_resize_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_resize_1/index_resize_req
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_resize_1/index_resize_ack
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_scale_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_scale_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_scale_1/scale_rename_req
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_index_scale_1/scale_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_final_index_sum_regn_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_final_index_sum_regn_Sample/req
      -- 
    ca_7169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2600_inst_ack_1, ack => convTransposeC_CP_6511_elements(40)); -- 
    req_7194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(40), ack => array_obj_ref_2606_index_offset_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_final_index_sum_regn_sample_complete
      -- CP-element group 41: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_final_index_sum_regn_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_final_index_sum_regn_Sample/ack
      -- 
    ack_7195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2606_index_offset_ack_0, ack => convTransposeC_CP_6511_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	92 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_offset_calculated
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_final_index_sum_regn_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_final_index_sum_regn_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_request/$entry
      -- CP-element group 42: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_request/req
      -- 
    ack_7200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2606_index_offset_ack_1, ack => convTransposeC_CP_6511_elements(42)); -- 
    req_7209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(42), ack => addr_of_2607_final_reg_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_request/$exit
      -- CP-element group 43: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_request/ack
      -- 
    ack_7210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2607_final_reg_ack_0, ack => convTransposeC_CP_6511_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	92 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (24) 
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_complete/ack
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_base_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_word_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_base_address_resized
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_base_addr_resize/$entry
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_base_addr_resize/$exit
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_base_addr_resize/base_resize_req
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_base_addr_resize/base_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_word_addrgen/$entry
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_word_addrgen/$exit
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_word_addrgen/root_register_req
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_word_addrgen/root_register_ack
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Sample/word_access_start/word_0/rr
      -- 
    ack_7215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2607_final_reg_ack_1, ack => convTransposeC_CP_6511_elements(44)); -- 
    rr_7248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(44), ack => ptr_deref_2611_load_0_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Sample/word_access_start/word_0/ra
      -- 
    ra_7249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2611_load_0_ack_0, ack => convTransposeC_CP_6511_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	92 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	53 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/ptr_deref_2611_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/ptr_deref_2611_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/ptr_deref_2611_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/ptr_deref_2611_Merge/merge_ack
      -- 
    ca_7260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2611_load_0_ack_1, ack => convTransposeC_CP_6511_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_Sample/ra
      -- 
    ra_7274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2631_inst_ack_0, ack => convTransposeC_CP_6511_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	92 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (16) 
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_resized_1
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_scaled_1
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_computed_1
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_resize_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_resize_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_resize_1/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_resize_1/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_scale_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_scale_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_scale_1/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_index_scale_1/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_final_index_sum_regn_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_final_index_sum_regn_Sample/req
      -- 
    ca_7279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2631_inst_ack_1, ack => convTransposeC_CP_6511_elements(48)); -- 
    req_7304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(48), ack => array_obj_ref_2637_index_offset_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_final_index_sum_regn_sample_complete
      -- CP-element group 49: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_final_index_sum_regn_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_final_index_sum_regn_Sample/ack
      -- 
    ack_7305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2637_index_offset_ack_0, ack => convTransposeC_CP_6511_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	92 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (11) 
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_request/req
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_request/$entry
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_offset_calculated
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_final_index_sum_regn_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_final_index_sum_regn_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_base_plus_offset/sum_rename_ack
      -- 
    ack_7310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2637_index_offset_ack_1, ack => convTransposeC_CP_6511_elements(50)); -- 
    req_7319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(50), ack => addr_of_2638_final_reg_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_request/ack
      -- CP-element group 51: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_request/$exit
      -- CP-element group 51: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_sample_completed_
      -- 
    ack_7320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2638_final_reg_ack_0, ack => convTransposeC_CP_6511_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	92 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (19) 
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_complete/ack
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_update_completed_
      -- 
    ack_7325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2638_final_reg_ack_1, ack => convTransposeC_CP_6511_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	46 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/word_access_start/word_0/rr
      -- CP-element group 53: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/ptr_deref_2641_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/ptr_deref_2641_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/ptr_deref_2641_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/ptr_deref_2641_Split/$entry
      -- 
    rr_7363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(53), ack => ptr_deref_2641_store_0_req_0); -- 
    convTransposeC_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(46) & convTransposeC_CP_6511_elements(52);
      gj_convTransposeC_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/word_access_start/word_0/ra
      -- CP-element group 54: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Sample/word_access_start/$exit
      -- 
    ra_7364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2641_store_0_ack_0, ack => convTransposeC_CP_6511_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	92 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Update/word_access_complete/$exit
      -- 
    ca_7375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2641_store_0_ack_1, ack => convTransposeC_CP_6511_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	92 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_sample_completed_
      -- 
    ra_7384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2647_inst_ack_0, ack => convTransposeC_CP_6511_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	92 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_Update/ca
      -- 
    ca_7389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2647_inst_ack_1, ack => convTransposeC_CP_6511_elements(57)); -- 
    -- CP-element group 58:  branch  join  transition  place  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659__exit__
      -- CP-element group 58: 	 branch_block_stmt_2284/if_stmt_2660__entry__
      -- CP-element group 58: 	 branch_block_stmt_2284/R_cmp_2661_place
      -- CP-element group 58: 	 branch_block_stmt_2284/if_stmt_2660_else_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2284/if_stmt_2660_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2284/if_stmt_2660_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_2284/if_stmt_2660_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_2284/if_stmt_2660_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_2284/if_stmt_2660_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/$exit
      -- 
    branch_req_7397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(58), ack => if_stmt_2660_branch_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(41) & convTransposeC_CP_6511_elements(49) & convTransposeC_CP_6511_elements(55) & convTransposeC_CP_6511_elements(57);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	87 
    -- CP-element group 59: 	88 
    -- CP-element group 59:  members (24) 
      -- CP-element group 59: 	 branch_block_stmt_2284/merge_stmt_2666__exit__
      -- CP-element group 59: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody
      -- CP-element group 59: 	 branch_block_stmt_2284/assign_stmt_2672__entry__
      -- CP-element group 59: 	 branch_block_stmt_2284/merge_stmt_2666_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_2284/assign_stmt_2672__exit__
      -- CP-element group 59: 	 branch_block_stmt_2284/whilex_xbody_ifx_xthen
      -- CP-element group 59: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/$entry
      -- CP-element group 59: 	 branch_block_stmt_2284/assign_stmt_2672/$entry
      -- CP-element group 59: 	 branch_block_stmt_2284/assign_stmt_2672/$exit
      -- CP-element group 59: 	 branch_block_stmt_2284/if_stmt_2660_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_2284/if_stmt_2660_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/$entry
      -- CP-element group 59: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_2284/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_2284/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_2284/merge_stmt_2666_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_2284/merge_stmt_2666_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_2284/merge_stmt_2666_PhiAck/dummy
      -- 
    if_choice_transition_7402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2660_branch_ack_1, ack => convTransposeC_CP_6511_elements(59)); -- 
    rr_7600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(59), ack => type_cast_2560_inst_req_0); -- 
    cr_7605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(59), ack => type_cast_2560_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	64 
    -- CP-element group 60: 	66 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (24) 
      -- CP-element group 60: 	 branch_block_stmt_2284/merge_stmt_2674_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_2284/merge_stmt_2674__exit__
      -- CP-element group 60: 	 branch_block_stmt_2284/whilex_xbody_ifx_xelse
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/$entry
      -- CP-element group 60: 	 branch_block_stmt_2284/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716__entry__
      -- CP-element group 60: 	 branch_block_stmt_2284/if_stmt_2660_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_2284/if_stmt_2660_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2284/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_2284/merge_stmt_2674_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_2284/merge_stmt_2674_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_2284/merge_stmt_2674_PhiAck/dummy
      -- 
    else_choice_transition_7406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2660_branch_ack_0, ack => convTransposeC_CP_6511_elements(60)); -- 
    cr_7455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(60), ack => type_cast_2710_inst_req_1); -- 
    cr_7441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(60), ack => type_cast_2693_inst_req_1); -- 
    cr_7427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(60), ack => type_cast_2684_inst_req_1); -- 
    rr_7422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(60), ack => type_cast_2684_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_Sample/$exit
      -- 
    ra_7423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2684_inst_ack_0, ack => convTransposeC_CP_6511_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2684_update_completed_
      -- 
    ca_7428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2684_inst_ack_1, ack => convTransposeC_CP_6511_elements(62)); -- 
    rr_7436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(62), ack => type_cast_2693_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_sample_completed_
      -- 
    ra_7437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2693_inst_ack_0, ack => convTransposeC_CP_6511_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	60 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2693_update_completed_
      -- 
    ca_7442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2693_inst_ack_1, ack => convTransposeC_CP_6511_elements(64)); -- 
    rr_7450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(64), ack => type_cast_2710_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_Sample/ra
      -- CP-element group 65: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_sample_completed_
      -- 
    ra_7451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2710_inst_ack_0, ack => convTransposeC_CP_6511_elements(65)); -- 
    -- CP-element group 66:  branch  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	60 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (13) 
      -- CP-element group 66: 	 branch_block_stmt_2284/R_cmp87_2718_place
      -- CP-element group 66: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716__exit__
      -- CP-element group 66: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/$exit
      -- CP-element group 66: 	 branch_block_stmt_2284/if_stmt_2717__entry__
      -- CP-element group 66: 	 branch_block_stmt_2284/if_stmt_2717_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2284/if_stmt_2717_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2284/if_stmt_2717_else_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2284/if_stmt_2717_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2284/if_stmt_2717_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2284/if_stmt_2717_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2284/assign_stmt_2680_to_assign_stmt_2716/type_cast_2710_update_completed_
      -- 
    ca_7456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2710_inst_ack_1, ack => convTransposeC_CP_6511_elements(66)); -- 
    branch_req_7464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(66), ack => if_stmt_2717_branch_req_0); -- 
    -- CP-element group 67:  merge  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (15) 
      -- CP-element group 67: 	 branch_block_stmt_2284/merge_stmt_2723__exit__
      -- CP-element group 67: 	 branch_block_stmt_2284/ifx_xelse_whilex_xend
      -- CP-element group 67: 	 branch_block_stmt_2284/assign_stmt_2727__entry__
      -- CP-element group 67: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_Sample/req
      -- CP-element group 67: 	 branch_block_stmt_2284/assign_stmt_2727/$entry
      -- CP-element group 67: 	 branch_block_stmt_2284/if_stmt_2717_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2284/if_stmt_2717_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_2284/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2284/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2284/merge_stmt_2723_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2284/merge_stmt_2723_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2284/merge_stmt_2723_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2284/merge_stmt_2723_PhiAck/dummy
      -- 
    if_choice_transition_7469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2717_branch_ack_1, ack => convTransposeC_CP_6511_elements(67)); -- 
    req_7486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(67), ack => WPIPE_Block2_done_2725_inst_req_0); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	77 
    -- CP-element group 68: 	79 
    -- CP-element group 68: 	80 
    -- CP-element group 68: 	76 
    -- CP-element group 68:  members (20) 
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/if_stmt_2717_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2284/if_stmt_2717_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/SplitProtocol/Update/$entry
      -- 
    else_choice_transition_7473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2717_branch_ack_0, ack => convTransposeC_CP_6511_elements(68)); -- 
    rr_7568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(68), ack => type_cast_2438_inst_req_0); -- 
    rr_7545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(68), ack => type_cast_2432_inst_req_0); -- 
    cr_7573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(68), ack => type_cast_2438_inst_req_1); -- 
    cr_7550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(68), ack => type_cast_2432_inst_req_1); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_Update/req
      -- CP-element group 69: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_Sample/ack
      -- CP-element group 69: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_update_start_
      -- CP-element group 69: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_sample_completed_
      -- 
    ack_7487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2725_inst_ack_0, ack => convTransposeC_CP_6511_elements(69)); -- 
    req_7491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(69), ack => WPIPE_Block2_done_2725_inst_req_1); -- 
    -- CP-element group 70:  transition  place  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (16) 
      -- CP-element group 70: 	 branch_block_stmt_2284/branch_block_stmt_2284__exit__
      -- CP-element group 70: 	 $exit
      -- CP-element group 70: 	 branch_block_stmt_2284/$exit
      -- CP-element group 70: 	 branch_block_stmt_2284/return__
      -- CP-element group 70: 	 branch_block_stmt_2284/merge_stmt_2729__exit__
      -- CP-element group 70: 	 branch_block_stmt_2284/assign_stmt_2727__exit__
      -- CP-element group 70: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2284/assign_stmt_2727/$exit
      -- CP-element group 70: 	 branch_block_stmt_2284/assign_stmt_2727/WPIPE_Block2_done_2725_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2284/return___PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2284/return___PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2284/merge_stmt_2729_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2284/merge_stmt_2729_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2284/merge_stmt_2729_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2284/merge_stmt_2729_PhiAck/dummy
      -- 
    ack_7492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2725_inst_ack_1, ack => convTransposeC_CP_6511_elements(70)); -- 
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	75 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2430_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/$exit
      -- CP-element group 71: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_req
      -- 
    phi_stmt_2426_req_7503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2426_req_7503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(71), ack => phi_stmt_2426_req_0); -- 
    -- Element group convTransposeC_CP_6511_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeC_CP_6511_elements(31), ack => convTransposeC_CP_6511_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	31 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Sample/$exit
      -- 
    ra_7520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2436_inst_ack_0, ack => convTransposeC_CP_6511_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	31 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Update/ca
      -- CP-element group 73: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/Update/$exit
      -- 
    ca_7525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2436_inst_ack_1, ack => convTransposeC_CP_6511_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/$exit
      -- CP-element group 74: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_req
      -- CP-element group 74: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2436/$exit
      -- CP-element group 74: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/$exit
      -- 
    phi_stmt_2433_req_7526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2433_req_7526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(74), ack => phi_stmt_2433_req_0); -- 
    convTransposeC_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(72) & convTransposeC_CP_6511_elements(73);
      gj_convTransposeC_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: 	71 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	83 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_2284/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(74) & convTransposeC_CP_6511_elements(71);
      gj_convTransposeC_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	68 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/SplitProtocol/Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/SplitProtocol/Sample/ra
      -- 
    ra_7546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2432_inst_ack_0, ack => convTransposeC_CP_6511_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	68 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/SplitProtocol/Update/ca
      -- CP-element group 77: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/SplitProtocol/Update/$exit
      -- 
    ca_7551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2432_inst_ack_1, ack => convTransposeC_CP_6511_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	82 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/type_cast_2432/$exit
      -- CP-element group 78: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/$exit
      -- CP-element group 78: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2426/phi_stmt_2426_req
      -- 
    phi_stmt_2426_req_7552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2426_req_7552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(78), ack => phi_stmt_2426_req_1); -- 
    convTransposeC_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(77) & convTransposeC_CP_6511_elements(76);
      gj_convTransposeC_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	68 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Sample/ra
      -- 
    ra_7569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2438_inst_ack_0, ack => convTransposeC_CP_6511_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	68 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Update/ca
      -- CP-element group 80: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/Update/$exit
      -- 
    ca_7574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2438_inst_ack_1, ack => convTransposeC_CP_6511_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_req
      -- CP-element group 81: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/type_cast_2438/$exit
      -- CP-element group 81: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/$exit
      -- CP-element group 81: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2433/phi_stmt_2433_sources/$exit
      -- 
    phi_stmt_2433_req_7575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2433_req_7575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(81), ack => phi_stmt_2433_req_1); -- 
    convTransposeC_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(79) & convTransposeC_CP_6511_elements(80);
      gj_convTransposeC_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2284/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(78) & convTransposeC_CP_6511_elements(81);
      gj_convTransposeC_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  merge  fork  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: 	75 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2284/merge_stmt_2425_PhiReqMerge
      -- CP-element group 83: 	 branch_block_stmt_2284/merge_stmt_2425_PhiAck/$entry
      -- 
    convTransposeC_CP_6511_elements(83) <= OrReduce(convTransposeC_CP_6511_elements(82) & convTransposeC_CP_6511_elements(75));
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2284/merge_stmt_2425_PhiAck/phi_stmt_2426_ack
      -- 
    phi_stmt_2426_ack_7580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2426_ack_0, ack => convTransposeC_CP_6511_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2284/merge_stmt_2425_PhiAck/phi_stmt_2433_ack
      -- 
    phi_stmt_2433_ack_7581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2433_ack_0, ack => convTransposeC_CP_6511_elements(85)); -- 
    -- CP-element group 86:  join  fork  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	34 
    -- CP-element group 86: 	35 
    -- CP-element group 86: 	32 
    -- CP-element group 86: 	33 
    -- CP-element group 86:  members (16) 
      -- CP-element group 86: 	 branch_block_stmt_2284/merge_stmt_2425__exit__
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551__entry__
      -- CP-element group 86: 	 branch_block_stmt_2284/merge_stmt_2425_PhiAck/$exit
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/$entry
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2443_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2284/assign_stmt_2444_to_assign_stmt_2551/type_cast_2448_Update/cr
      -- 
    rr_7118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(86), ack => type_cast_2443_inst_req_0); -- 
    cr_7123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(86), ack => type_cast_2443_inst_req_1); -- 
    rr_7132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(86), ack => type_cast_2448_inst_req_0); -- 
    cr_7137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(86), ack => type_cast_2448_inst_req_1); -- 
    convTransposeC_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(84) & convTransposeC_CP_6511_elements(85);
      gj_convTransposeC_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	59 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/SplitProtocol/Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/SplitProtocol/Sample/$exit
      -- 
    ra_7601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2560_inst_ack_0, ack => convTransposeC_CP_6511_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	59 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/SplitProtocol/Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/SplitProtocol/Update/ca
      -- 
    ca_7606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2560_inst_ack_1, ack => convTransposeC_CP_6511_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/$exit
      -- CP-element group 89: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/$exit
      -- CP-element group 89: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 89: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2560/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_2284/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_req
      -- 
    phi_stmt_2554_req_7607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2554_req_7607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(89), ack => phi_stmt_2554_req_1); -- 
    convTransposeC_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(87) & convTransposeC_CP_6511_elements(88);
      gj_convTransposeC_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  output  delay-element  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	36 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2284/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_2284/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2554/$exit
      -- CP-element group 90: 	 branch_block_stmt_2284/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2284/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_sources/type_cast_2558_konst_delay_trans
      -- CP-element group 90: 	 branch_block_stmt_2284/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2554/phi_stmt_2554_req
      -- 
    phi_stmt_2554_req_7618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2554_req_7618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(90), ack => phi_stmt_2554_req_0); -- 
    -- Element group convTransposeC_CP_6511_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => convTransposeC_CP_6511_elements(36), ack => convTransposeC_CP_6511_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  merge  transition  place  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2284/merge_stmt_2553_PhiReqMerge
      -- CP-element group 91: 	 branch_block_stmt_2284/merge_stmt_2553_PhiAck/$entry
      -- 
    convTransposeC_CP_6511_elements(91) <= OrReduce(convTransposeC_CP_6511_elements(90) & convTransposeC_CP_6511_elements(89));
    -- CP-element group 92:  fork  transition  place  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	40 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	38 
    -- CP-element group 92: 	42 
    -- CP-element group 92: 	44 
    -- CP-element group 92: 	46 
    -- CP-element group 92: 	48 
    -- CP-element group 92: 	50 
    -- CP-element group 92: 	52 
    -- CP-element group 92: 	55 
    -- CP-element group 92: 	56 
    -- CP-element group 92: 	57 
    -- CP-element group 92:  members (45) 
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659__entry__
      -- CP-element group 92: 	 branch_block_stmt_2284/merge_stmt_2553__exit__
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2647_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2641_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2570_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2600_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2606_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2607_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/ptr_deref_2611_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/type_cast_2631_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/addr_of_2638_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2284/assign_stmt_2567_to_assign_stmt_2659/array_obj_ref_2637_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2284/merge_stmt_2553_PhiAck/$exit
      -- CP-element group 92: 	 branch_block_stmt_2284/merge_stmt_2553_PhiAck/phi_stmt_2554_ack
      -- 
    phi_stmt_2554_ack_7623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2554_ack_0, ack => convTransposeC_CP_6511_elements(92)); -- 
    cr_7388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2647_inst_req_1); -- 
    rr_7383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2647_inst_req_0); -- 
    cr_7374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => ptr_deref_2641_store_0_req_1); -- 
    req_7324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => addr_of_2638_final_reg_req_1); -- 
    rr_7149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2570_inst_req_0); -- 
    cr_7154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2570_inst_req_1); -- 
    cr_7168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2600_inst_req_1); -- 
    req_7199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => array_obj_ref_2606_index_offset_req_1); -- 
    req_7214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => addr_of_2607_final_reg_req_1); -- 
    cr_7259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => ptr_deref_2611_load_0_req_1); -- 
    cr_7278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2631_inst_req_1); -- 
    req_7309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => array_obj_ref_2637_index_offset_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2513_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2534_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2594_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2625_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2362_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2362_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom62_2636_resized : std_logic_vector(13 downto 0);
    signal R_idxprom62_2636_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2605_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2605_scaled : std_logic_vector(13 downto 0);
    signal add18_2576 : std_logic_vector(31 downto 0);
    signal add26_2474 : std_logic_vector(31 downto 0);
    signal add37_2489 : std_logic_vector(31 downto 0);
    signal add52_2546 : std_logic_vector(31 downto 0);
    signal add54_2581 : std_logic_vector(31 downto 0);
    signal add67_2654 : std_logic_vector(31 downto 0);
    signal add_2459 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2606_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2606_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2606_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2606_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2606_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2606_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2637_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2637_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2637_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2637_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2637_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2637_root_address : std_logic_vector(13 downto 0);
    signal arrayidx63_2639 : std_logic_vector(31 downto 0);
    signal arrayidx_2608 : std_logic_vector(31 downto 0);
    signal call_2287 : std_logic_vector(15 downto 0);
    signal cmp79_2690 : std_logic_vector(0 downto 0);
    signal cmp87_2716 : std_logic_vector(0 downto 0);
    signal cmp_2659 : std_logic_vector(0 downto 0);
    signal conv10100_2571 : std_logic_vector(31 downto 0);
    signal conv13_2444 : std_logic_vector(31 downto 0);
    signal conv16_2449 : std_logic_vector(31 downto 0);
    signal conv23_2348 : std_logic_vector(31 downto 0);
    signal conv28_2367 : std_logic_vector(31 downto 0);
    signal conv34_2381 : std_logic_vector(31 downto 0);
    signal conv47_2515 : std_logic_vector(31 downto 0);
    signal conv50_2536 : std_logic_vector(31 downto 0);
    signal conv66_2648 : std_logic_vector(31 downto 0);
    signal conv76_2685 : std_logic_vector(31 downto 0);
    signal conv85_2711 : std_logic_vector(31 downto 0);
    signal conv_2310 : std_logic_vector(15 downto 0);
    signal div78_2423 : std_logic_vector(31 downto 0);
    signal div_2306 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2413 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2296 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2318 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2330 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2340 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2356 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2373 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2389 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2401 : std_logic_vector(31 downto 0);
    signal idxprom62_2632 : std_logic_vector(63 downto 0);
    signal idxprom_2601 : std_logic_vector(63 downto 0);
    signal inc83_2694 : std_logic_vector(15 downto 0);
    signal inc83x_xinput_dim0x_x2_2699 : std_logic_vector(15 downto 0);
    signal inc_2680 : std_logic_vector(15 downto 0);
    signal indvar_2554 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2672 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2433 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2426 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2706 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2567 : std_logic_vector(15 downto 0);
    signal mul17_2464 : std_logic_vector(31 downto 0);
    signal mul24_2469 : std_logic_vector(31 downto 0);
    signal mul35_2484 : std_logic_vector(31 downto 0);
    signal mul51_2541 : std_logic_vector(31 downto 0);
    signal mul53_2551 : std_logic_vector(31 downto 0);
    signal mul_2454 : std_logic_vector(31 downto 0);
    signal ptr_deref_2299_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2299_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2299_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2299_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2299_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2321_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2321_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2321_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2321_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2321_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2333_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2333_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2333_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2333_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2333_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2343_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2343_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2343_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2343_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2343_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2359_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2359_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2359_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2359_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2359_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2376_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2376_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2376_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2376_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2376_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2392_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2392_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2392_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2392_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2392_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2404_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2404_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2404_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2404_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2404_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2416_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2416_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2416_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2416_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2416_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2611_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2611_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2611_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2611_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2611_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2641_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2641_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2641_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2641_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2641_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2641_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext101_2527 : std_logic_vector(31 downto 0);
    signal sext103_2587 : std_logic_vector(31 downto 0);
    signal sext104_2618 : std_logic_vector(31 downto 0);
    signal sext_2506 : std_logic_vector(31 downto 0);
    signal shr61_2627 : std_logic_vector(31 downto 0);
    signal shr_2596 : std_logic_vector(31 downto 0);
    signal sub29_2521 : std_logic_vector(31 downto 0);
    signal sub40_2494 : std_logic_vector(31 downto 0);
    signal sub41_2500 : std_logic_vector(31 downto 0);
    signal sub_2479 : std_logic_vector(31 downto 0);
    signal tmp11_2322 : std_logic_vector(31 downto 0);
    signal tmp14_2334 : std_logic_vector(31 downto 0);
    signal tmp22_2344 : std_logic_vector(15 downto 0);
    signal tmp25_2360 : std_logic_vector(31 downto 0);
    signal tmp27_2363 : std_logic_vector(15 downto 0);
    signal tmp33_2377 : std_logic_vector(15 downto 0);
    signal tmp36_2393 : std_logic_vector(31 downto 0);
    signal tmp45_2405 : std_logic_vector(31 downto 0);
    signal tmp48_2417 : std_logic_vector(31 downto 0);
    signal tmp58_2612 : std_logic_vector(63 downto 0);
    signal tmp_2300 : std_logic_vector(31 downto 0);
    signal type_cast_2304_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2421_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2430_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2432_wire : std_logic_vector(15 downto 0);
    signal type_cast_2436_wire : std_logic_vector(15 downto 0);
    signal type_cast_2438_wire : std_logic_vector(15 downto 0);
    signal type_cast_2442_wire : std_logic_vector(31 downto 0);
    signal type_cast_2447_wire : std_logic_vector(31 downto 0);
    signal type_cast_2498_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2504_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2509_wire : std_logic_vector(31 downto 0);
    signal type_cast_2512_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2519_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2525_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2530_wire : std_logic_vector(31 downto 0);
    signal type_cast_2533_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2558_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2560_wire : std_logic_vector(15 downto 0);
    signal type_cast_2565_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2585_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2590_wire : std_logic_vector(31 downto 0);
    signal type_cast_2593_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2599_wire : std_logic_vector(63 downto 0);
    signal type_cast_2616_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2621_wire : std_logic_vector(31 downto 0);
    signal type_cast_2624_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2630_wire : std_logic_vector(63 downto 0);
    signal type_cast_2646_wire : std_logic_vector(31 downto 0);
    signal type_cast_2652_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2670_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2678_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2683_wire : std_logic_vector(31 downto 0);
    signal type_cast_2703_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2709_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2362_word_address_0 <= "0";
    array_obj_ref_2606_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2606_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2606_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2606_resized_base_address <= "00000000000000";
    array_obj_ref_2637_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2637_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2637_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2637_resized_base_address <= "00000000000000";
    iNsTr_10_2413 <= "00000000000000000000000000000011";
    iNsTr_2_2296 <= "00000000000000000000000000000010";
    iNsTr_3_2318 <= "00000000000000000000000000000100";
    iNsTr_4_2330 <= "00000000000000000000000000000011";
    iNsTr_5_2340 <= "00000000000000000000000000000000";
    iNsTr_6_2356 <= "00000000000000000000000000000011";
    iNsTr_7_2373 <= "00000000000000000000000000000001";
    iNsTr_8_2389 <= "00000000000000000000000000000100";
    iNsTr_9_2401 <= "00000000000000000000000000000100";
    ptr_deref_2299_word_offset_0 <= "0000000";
    ptr_deref_2321_word_offset_0 <= "0000000";
    ptr_deref_2333_word_offset_0 <= "0000000";
    ptr_deref_2343_word_offset_0 <= "0";
    ptr_deref_2359_word_offset_0 <= "0000000";
    ptr_deref_2376_word_offset_0 <= "0";
    ptr_deref_2392_word_offset_0 <= "0000000";
    ptr_deref_2404_word_offset_0 <= "0000000";
    ptr_deref_2416_word_offset_0 <= "0000000";
    ptr_deref_2611_word_offset_0 <= "00000000000000";
    ptr_deref_2641_word_offset_0 <= "00000000000000";
    type_cast_2304_wire_constant <= "00000000000000000000000000000001";
    type_cast_2421_wire_constant <= "00000000000000000000000000000001";
    type_cast_2430_wire_constant <= "0000000000000000";
    type_cast_2498_wire_constant <= "00000000000000000000000000010000";
    type_cast_2504_wire_constant <= "11111111111111110000000000000000";
    type_cast_2512_wire_constant <= "00000000000000000000000000010000";
    type_cast_2519_wire_constant <= "00000000000000000000000000010000";
    type_cast_2525_wire_constant <= "11111111111111110000000000000000";
    type_cast_2533_wire_constant <= "00000000000000000000000000010000";
    type_cast_2558_wire_constant <= "0000000000000000";
    type_cast_2565_wire_constant <= "0000000000000100";
    type_cast_2585_wire_constant <= "00000000000000000000000000010000";
    type_cast_2593_wire_constant <= "00000000000000000000000000010010";
    type_cast_2616_wire_constant <= "00000000000000000000000000010000";
    type_cast_2624_wire_constant <= "00000000000000000000000000010010";
    type_cast_2652_wire_constant <= "00000000000000000000000000000100";
    type_cast_2670_wire_constant <= "0000000000000001";
    type_cast_2678_wire_constant <= "0000000000000001";
    type_cast_2703_wire_constant <= "0000000000000000";
    phi_stmt_2426: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2430_wire_constant & type_cast_2432_wire;
      req <= phi_stmt_2426_req_0 & phi_stmt_2426_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2426",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2426_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2426,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2426
    phi_stmt_2433: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2436_wire & type_cast_2438_wire;
      req <= phi_stmt_2433_req_0 & phi_stmt_2433_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2433",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2433_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2433,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2433
    phi_stmt_2554: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2558_wire_constant & type_cast_2560_wire;
      req <= phi_stmt_2554_req_0 & phi_stmt_2554_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2554",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2554_ack_0,
          idata => idata,
          odata => indvar_2554,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2554
    -- flow-through select operator MUX_2705_inst
    input_dim1x_x2_2706 <= type_cast_2703_wire_constant when (cmp79_2690(0) /=  '0') else inc_2680;
    addr_of_2607_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2607_final_reg_req_0;
      addr_of_2607_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2607_final_reg_req_1;
      addr_of_2607_final_reg_ack_1<= rack(0);
      addr_of_2607_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2607_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2606_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2608,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2638_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2638_final_reg_req_0;
      addr_of_2638_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2638_final_reg_req_1;
      addr_of_2638_final_reg_ack_1<= rack(0);
      addr_of_2638_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2638_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2637_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx63_2639,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2309_inst_req_0;
      type_cast_2309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2309_inst_req_1;
      type_cast_2309_inst_ack_1<= rack(0);
      type_cast_2309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2306,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2310,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2347_inst_req_0;
      type_cast_2347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2347_inst_req_1;
      type_cast_2347_inst_ack_1<= rack(0);
      type_cast_2347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp22_2344,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_2348,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2366_inst_req_0;
      type_cast_2366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2366_inst_req_1;
      type_cast_2366_inst_ack_1<= rack(0);
      type_cast_2366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp27_2363,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28_2367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2380_inst_req_0;
      type_cast_2380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2380_inst_req_1;
      type_cast_2380_inst_ack_1<= rack(0);
      type_cast_2380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp33_2377,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34_2381,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2432_inst_req_0;
      type_cast_2432_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2432_inst_req_1;
      type_cast_2432_inst_ack_1<= rack(0);
      type_cast_2432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2706,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2432_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2436_inst_req_0;
      type_cast_2436_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2436_inst_req_1;
      type_cast_2436_inst_ack_1<= rack(0);
      type_cast_2436_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2310,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2436_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2438_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2438_inst_req_0;
      type_cast_2438_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2438_inst_req_1;
      type_cast_2438_inst_ack_1<= rack(0);
      type_cast_2438_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2438_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc83x_xinput_dim0x_x2_2699,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2438_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2443_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2443_inst_req_0;
      type_cast_2443_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2443_inst_req_1;
      type_cast_2443_inst_ack_1<= rack(0);
      type_cast_2443_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2443_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2442_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_2444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2448_inst_req_0;
      type_cast_2448_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2448_inst_req_1;
      type_cast_2448_inst_ack_1<= rack(0);
      type_cast_2448_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2448_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2447_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_2449,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2509_inst
    process(sext_2506) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2506(31 downto 0);
      type_cast_2509_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2514_inst
    process(ASHR_i32_i32_2513_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2513_wire(31 downto 0);
      conv47_2515 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2530_inst
    process(sext101_2527) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext101_2527(31 downto 0);
      type_cast_2530_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2535_inst
    process(ASHR_i32_i32_2534_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2534_wire(31 downto 0);
      conv50_2536 <= tmp_var; -- 
    end process;
    type_cast_2560_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2560_inst_req_0;
      type_cast_2560_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2560_inst_req_1;
      type_cast_2560_inst_ack_1<= rack(0);
      type_cast_2560_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2560_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2672,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2560_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2570_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2570_inst_req_0;
      type_cast_2570_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2570_inst_req_1;
      type_cast_2570_inst_ack_1<= rack(0);
      type_cast_2570_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2570_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2567,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10100_2571,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2590_inst
    process(sext103_2587) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext103_2587(31 downto 0);
      type_cast_2590_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2595_inst
    process(ASHR_i32_i32_2594_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2594_wire(31 downto 0);
      shr_2596 <= tmp_var; -- 
    end process;
    type_cast_2600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2600_inst_req_0;
      type_cast_2600_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2600_inst_req_1;
      type_cast_2600_inst_ack_1<= rack(0);
      type_cast_2600_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2600_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2599_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2601,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2621_inst
    process(sext104_2618) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext104_2618(31 downto 0);
      type_cast_2621_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2626_inst
    process(ASHR_i32_i32_2625_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2625_wire(31 downto 0);
      shr61_2627 <= tmp_var; -- 
    end process;
    type_cast_2631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2631_inst_req_0;
      type_cast_2631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2631_inst_req_1;
      type_cast_2631_inst_ack_1<= rack(0);
      type_cast_2631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2630_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom62_2632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2647_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2647_inst_req_0;
      type_cast_2647_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2647_inst_req_1;
      type_cast_2647_inst_ack_1<= rack(0);
      type_cast_2647_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2647_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2646_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_2648,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2684_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2684_inst_req_0;
      type_cast_2684_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2684_inst_req_1;
      type_cast_2684_inst_ack_1<= rack(0);
      type_cast_2684_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2684_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2683_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_2685,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2693_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2693_inst_req_0;
      type_cast_2693_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2693_inst_req_1;
      type_cast_2693_inst_ack_1<= rack(0);
      type_cast_2693_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2693_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp79_2690,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc83_2694,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2710_inst_req_0;
      type_cast_2710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2710_inst_req_1;
      type_cast_2710_inst_ack_1<= rack(0);
      type_cast_2710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2709_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_2711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2362_gather_scatter
    process(LOAD_padding_2362_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2362_data_0;
      ov(15 downto 0) := iv;
      tmp27_2363 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2606_index_1_rename
    process(R_idxprom_2605_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2605_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2605_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2606_index_1_resize
    process(idxprom_2601) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2601;
      ov := iv(13 downto 0);
      R_idxprom_2605_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2606_root_address_inst
    process(array_obj_ref_2606_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2606_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2606_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2637_index_1_rename
    process(R_idxprom62_2636_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom62_2636_resized;
      ov(13 downto 0) := iv;
      R_idxprom62_2636_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2637_index_1_resize
    process(idxprom62_2632) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom62_2632;
      ov := iv(13 downto 0);
      R_idxprom62_2636_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2637_root_address_inst
    process(array_obj_ref_2637_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2637_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2637_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2299_addr_0
    process(ptr_deref_2299_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2299_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2299_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2299_base_resize
    process(iNsTr_2_2296) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2296;
      ov := iv(6 downto 0);
      ptr_deref_2299_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2299_gather_scatter
    process(ptr_deref_2299_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2299_data_0;
      ov(31 downto 0) := iv;
      tmp_2300 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2299_root_address_inst
    process(ptr_deref_2299_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2299_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2299_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2321_addr_0
    process(ptr_deref_2321_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2321_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2321_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2321_base_resize
    process(iNsTr_3_2318) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2318;
      ov := iv(6 downto 0);
      ptr_deref_2321_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2321_gather_scatter
    process(ptr_deref_2321_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2321_data_0;
      ov(31 downto 0) := iv;
      tmp11_2322 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2321_root_address_inst
    process(ptr_deref_2321_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2321_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2321_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2333_addr_0
    process(ptr_deref_2333_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2333_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2333_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2333_base_resize
    process(iNsTr_4_2330) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2330;
      ov := iv(6 downto 0);
      ptr_deref_2333_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2333_gather_scatter
    process(ptr_deref_2333_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2333_data_0;
      ov(31 downto 0) := iv;
      tmp14_2334 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2333_root_address_inst
    process(ptr_deref_2333_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2333_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2333_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2343_addr_0
    process(ptr_deref_2343_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2343_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2343_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2343_base_resize
    process(iNsTr_5_2340) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2340;
      ov := iv(0 downto 0);
      ptr_deref_2343_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2343_gather_scatter
    process(ptr_deref_2343_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2343_data_0;
      ov(15 downto 0) := iv;
      tmp22_2344 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2343_root_address_inst
    process(ptr_deref_2343_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2343_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2343_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2359_addr_0
    process(ptr_deref_2359_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2359_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2359_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2359_base_resize
    process(iNsTr_6_2356) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2356;
      ov := iv(6 downto 0);
      ptr_deref_2359_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2359_gather_scatter
    process(ptr_deref_2359_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2359_data_0;
      ov(31 downto 0) := iv;
      tmp25_2360 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2359_root_address_inst
    process(ptr_deref_2359_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2359_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2359_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2376_addr_0
    process(ptr_deref_2376_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2376_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2376_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2376_base_resize
    process(iNsTr_7_2373) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2373;
      ov := iv(0 downto 0);
      ptr_deref_2376_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2376_gather_scatter
    process(ptr_deref_2376_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2376_data_0;
      ov(15 downto 0) := iv;
      tmp33_2377 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2376_root_address_inst
    process(ptr_deref_2376_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2376_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2376_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2392_addr_0
    process(ptr_deref_2392_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2392_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2392_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2392_base_resize
    process(iNsTr_8_2389) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2389;
      ov := iv(6 downto 0);
      ptr_deref_2392_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2392_gather_scatter
    process(ptr_deref_2392_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2392_data_0;
      ov(31 downto 0) := iv;
      tmp36_2393 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2392_root_address_inst
    process(ptr_deref_2392_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2392_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2392_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2404_addr_0
    process(ptr_deref_2404_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2404_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2404_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2404_base_resize
    process(iNsTr_9_2401) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2401;
      ov := iv(6 downto 0);
      ptr_deref_2404_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2404_gather_scatter
    process(ptr_deref_2404_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2404_data_0;
      ov(31 downto 0) := iv;
      tmp45_2405 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2404_root_address_inst
    process(ptr_deref_2404_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2404_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2404_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2416_addr_0
    process(ptr_deref_2416_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2416_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2416_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2416_base_resize
    process(iNsTr_10_2413) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2413;
      ov := iv(6 downto 0);
      ptr_deref_2416_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2416_gather_scatter
    process(ptr_deref_2416_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2416_data_0;
      ov(31 downto 0) := iv;
      tmp48_2417 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2416_root_address_inst
    process(ptr_deref_2416_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2416_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2416_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2611_addr_0
    process(ptr_deref_2611_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2611_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2611_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2611_base_resize
    process(arrayidx_2608) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2608;
      ov := iv(13 downto 0);
      ptr_deref_2611_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2611_gather_scatter
    process(ptr_deref_2611_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2611_data_0;
      ov(63 downto 0) := iv;
      tmp58_2612 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2611_root_address_inst
    process(ptr_deref_2611_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2611_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2611_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2641_addr_0
    process(ptr_deref_2641_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2641_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2641_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2641_base_resize
    process(arrayidx63_2639) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx63_2639;
      ov := iv(13 downto 0);
      ptr_deref_2641_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2641_gather_scatter
    process(tmp58_2612) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp58_2612;
      ov(63 downto 0) := iv;
      ptr_deref_2641_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2641_root_address_inst
    process(ptr_deref_2641_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2641_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2641_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2660_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2659;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2660_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2660_branch_req_0,
          ack0 => if_stmt_2660_branch_ack_0,
          ack1 => if_stmt_2660_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2717_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp87_2716;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2717_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2717_branch_req_0,
          ack0 => if_stmt_2717_branch_ack_0,
          ack1 => if_stmt_2717_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2671_inst
    process(indvar_2554) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2554, type_cast_2670_wire_constant, tmp_var);
      indvarx_xnext_2672 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2679_inst
    process(input_dim1x_x1x_xph_2426) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2426, type_cast_2678_wire_constant, tmp_var);
      inc_2680 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2698_inst
    process(inc83_2694, input_dim0x_x2x_xph_2433) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc83_2694, input_dim0x_x2x_xph_2433, tmp_var);
      inc83x_xinput_dim0x_x2_2699 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2458_inst
    process(mul_2454, conv13_2444) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2454, conv13_2444, tmp_var);
      add_2459 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2473_inst
    process(mul24_2469, tmp25_2360) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul24_2469, tmp25_2360, tmp_var);
      add26_2474 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2488_inst
    process(mul35_2484, tmp36_2393) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul35_2484, tmp36_2393, tmp_var);
      add37_2489 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2505_inst
    process(sub41_2500) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub41_2500, type_cast_2504_wire_constant, tmp_var);
      sext_2506 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2526_inst
    process(sub29_2521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub29_2521, type_cast_2525_wire_constant, tmp_var);
      sext101_2527 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2545_inst
    process(conv47_2515, mul51_2541) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv47_2515, mul51_2541, tmp_var);
      add52_2546 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2575_inst
    process(mul17_2464, conv10100_2571) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul17_2464, conv10100_2571, tmp_var);
      add18_2576 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2580_inst
    process(mul53_2551, conv10100_2571) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul53_2551, conv10100_2571, tmp_var);
      add54_2581 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2653_inst
    process(conv66_2648) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv66_2648, type_cast_2652_wire_constant, tmp_var);
      add67_2654 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2513_inst
    process(type_cast_2509_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2509_wire, type_cast_2512_wire_constant, tmp_var);
      ASHR_i32_i32_2513_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2534_inst
    process(type_cast_2530_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2530_wire, type_cast_2533_wire_constant, tmp_var);
      ASHR_i32_i32_2534_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2594_inst
    process(type_cast_2590_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2590_wire, type_cast_2593_wire_constant, tmp_var);
      ASHR_i32_i32_2594_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2625_inst
    process(type_cast_2621_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2621_wire, type_cast_2624_wire_constant, tmp_var);
      ASHR_i32_i32_2625_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2689_inst
    process(conv76_2685, div78_2423) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv76_2685, div78_2423, tmp_var);
      cmp79_2690 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2715_inst
    process(conv85_2711, tmp_2300) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv85_2711, tmp_2300, tmp_var);
      cmp87_2716 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2305_inst
    process(tmp_2300) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2300, type_cast_2304_wire_constant, tmp_var);
      div_2306 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2422_inst
    process(tmp14_2334) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_2334, type_cast_2421_wire_constant, tmp_var);
      div78_2423 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2566_inst
    process(indvar_2554) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2554, type_cast_2565_wire_constant, tmp_var);
      input_dim2x_x1_2567 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2453_inst
    process(tmp14_2334, conv16_2449) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_2334, conv16_2449, tmp_var);
      mul_2454 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2463_inst
    process(add_2459, tmp11_2322) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2459, tmp11_2322, tmp_var);
      mul17_2464 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2468_inst
    process(conv23_2348, conv16_2449) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv23_2348, conv16_2449, tmp_var);
      mul24_2469 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2483_inst
    process(conv34_2381, conv13_2444) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv34_2381, conv13_2444, tmp_var);
      mul35_2484 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2540_inst
    process(tmp48_2417, conv50_2536) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_2417, conv50_2536, tmp_var);
      mul51_2541 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2550_inst
    process(add52_2546, tmp45_2405) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add52_2546, tmp45_2405, tmp_var);
      mul53_2551 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2499_inst
    process(sub40_2494) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub40_2494, type_cast_2498_wire_constant, tmp_var);
      sub41_2500 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2520_inst
    process(sub_2479) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2479, type_cast_2519_wire_constant, tmp_var);
      sub29_2521 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2586_inst
    process(add18_2576) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add18_2576, type_cast_2585_wire_constant, tmp_var);
      sext103_2587 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2617_inst
    process(add54_2581) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add54_2581, type_cast_2616_wire_constant, tmp_var);
      sext104_2618 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2478_inst
    process(add26_2474, conv28_2367) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add26_2474, conv28_2367, tmp_var);
      sub_2479 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2493_inst
    process(add37_2489, conv28_2367) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add37_2489, conv28_2367, tmp_var);
      sub40_2494 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2658_inst
    process(add67_2654, tmp11_2322) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add67_2654, tmp11_2322, tmp_var);
      cmp_2659 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_2606_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2605_scaled;
      array_obj_ref_2606_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2606_index_offset_req_0;
      array_obj_ref_2606_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2606_index_offset_req_1;
      array_obj_ref_2606_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_2637_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom62_2636_scaled;
      array_obj_ref_2637_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2637_index_offset_req_0;
      array_obj_ref_2637_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2637_index_offset_req_1;
      array_obj_ref_2637_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- unary operator type_cast_2442_inst
    process(input_dim1x_x1x_xph_2426) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_2426, tmp_var);
      type_cast_2442_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2447_inst
    process(input_dim0x_x2x_xph_2433) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_2433, tmp_var);
      type_cast_2447_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2599_inst
    process(shr_2596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2596, tmp_var);
      type_cast_2599_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2630_inst
    process(shr61_2627) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr61_2627, tmp_var);
      type_cast_2630_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2646_inst
    process(input_dim2x_x1_2567) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2567, tmp_var);
      type_cast_2646_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2683_inst
    process(inc_2680) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2680, tmp_var);
      type_cast_2683_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2709_inst
    process(inc83x_xinput_dim0x_x2_2699) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc83x_xinput_dim0x_x2_2699, tmp_var);
      type_cast_2709_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2362_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2362_load_0_req_0;
      LOAD_padding_2362_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2362_load_0_req_1;
      LOAD_padding_2362_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2362_word_address_0;
      LOAD_padding_2362_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2299_load_0 ptr_deref_2321_load_0 ptr_deref_2333_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2299_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2321_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2333_load_0_req_0;
      ptr_deref_2299_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2321_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2333_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2299_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2321_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2333_load_0_req_1;
      ptr_deref_2299_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2321_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2333_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2299_word_address_0 & ptr_deref_2321_word_address_0 & ptr_deref_2333_word_address_0;
      ptr_deref_2299_data_0 <= data_out(95 downto 64);
      ptr_deref_2321_data_0 <= data_out(63 downto 32);
      ptr_deref_2333_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2343_load_0 ptr_deref_2376_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2343_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2376_load_0_req_0;
      ptr_deref_2343_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2376_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2343_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2376_load_0_req_1;
      ptr_deref_2343_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2376_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2343_word_address_0 & ptr_deref_2376_word_address_0;
      ptr_deref_2343_data_0 <= data_out(31 downto 16);
      ptr_deref_2376_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2359_load_0 ptr_deref_2392_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2359_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2392_load_0_req_0;
      ptr_deref_2359_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2392_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2359_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2392_load_0_req_1;
      ptr_deref_2359_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2392_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2359_word_address_0 & ptr_deref_2392_word_address_0;
      ptr_deref_2359_data_0 <= data_out(63 downto 32);
      ptr_deref_2392_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2404_load_0 ptr_deref_2416_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2404_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2416_load_0_req_0;
      ptr_deref_2404_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2416_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2404_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2416_load_0_req_1;
      ptr_deref_2404_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2416_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2404_word_address_0 & ptr_deref_2416_word_address_0;
      ptr_deref_2404_data_0 <= data_out(63 downto 32);
      ptr_deref_2416_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2611_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2611_load_0_req_0;
      ptr_deref_2611_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2611_load_0_req_1;
      ptr_deref_2611_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2611_word_address_0;
      ptr_deref_2611_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2641_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2641_store_0_req_0;
      ptr_deref_2641_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2641_store_0_req_1;
      ptr_deref_2641_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2641_word_address_0;
      data_in <= ptr_deref_2641_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2286_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_start_2286_inst_req_0;
      RPIPE_Block2_start_2286_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_start_2286_inst_req_1;
      RPIPE_Block2_start_2286_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2287 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2725_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2725_inst_req_0;
      WPIPE_Block2_done_2725_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2725_inst_req_1;
      WPIPE_Block2_done_2725_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2287;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_7664_start: Boolean;
  signal convTransposeD_CP_7664_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2839_inst_ack_1 : boolean;
  signal type_cast_2839_inst_req_1 : boolean;
  signal ptr_deref_2863_load_0_ack_1 : boolean;
  signal ptr_deref_2875_load_0_ack_0 : boolean;
  signal ptr_deref_2875_load_0_req_0 : boolean;
  signal type_cast_2806_inst_ack_1 : boolean;
  signal type_cast_2806_inst_req_1 : boolean;
  signal LOAD_padding_2821_load_0_req_0 : boolean;
  signal LOAD_padding_2821_load_0_ack_0 : boolean;
  signal type_cast_2895_inst_ack_1 : boolean;
  signal type_cast_2900_inst_req_0 : boolean;
  signal type_cast_2895_inst_req_0 : boolean;
  signal type_cast_2895_inst_ack_0 : boolean;
  signal type_cast_2839_inst_ack_0 : boolean;
  signal ptr_deref_2851_load_0_ack_0 : boolean;
  signal type_cast_2900_inst_ack_0 : boolean;
  signal type_cast_2839_inst_req_0 : boolean;
  signal type_cast_2895_inst_req_1 : boolean;
  signal ptr_deref_2875_load_0_req_1 : boolean;
  signal ptr_deref_2875_load_0_ack_1 : boolean;
  signal type_cast_2900_inst_req_1 : boolean;
  signal ptr_deref_2863_load_0_req_0 : boolean;
  signal LOAD_padding_2821_load_0_req_1 : boolean;
  signal LOAD_padding_2821_load_0_ack_1 : boolean;
  signal type_cast_3022_inst_ack_0 : boolean;
  signal ptr_deref_2863_load_0_req_1 : boolean;
  signal type_cast_3022_inst_req_0 : boolean;
  signal type_cast_2900_inst_ack_1 : boolean;
  signal ptr_deref_2863_load_0_ack_0 : boolean;
  signal type_cast_2806_inst_ack_0 : boolean;
  signal type_cast_2806_inst_req_0 : boolean;
  signal ptr_deref_2818_load_0_ack_0 : boolean;
  signal RPIPE_Block3_start_2735_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2735_inst_ack_0 : boolean;
  signal ptr_deref_2818_load_0_req_0 : boolean;
  signal RPIPE_Block3_start_2735_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2735_inst_ack_1 : boolean;
  signal ptr_deref_2851_load_0_req_0 : boolean;
  signal ptr_deref_2748_load_0_req_0 : boolean;
  signal ptr_deref_2748_load_0_ack_0 : boolean;
  signal ptr_deref_2748_load_0_req_1 : boolean;
  signal ptr_deref_2748_load_0_ack_1 : boolean;
  signal type_cast_2825_inst_ack_1 : boolean;
  signal type_cast_2825_inst_req_1 : boolean;
  signal type_cast_2758_inst_req_0 : boolean;
  signal type_cast_2758_inst_ack_0 : boolean;
  signal type_cast_2758_inst_req_1 : boolean;
  signal type_cast_2758_inst_ack_1 : boolean;
  signal ptr_deref_2835_load_0_ack_1 : boolean;
  signal ptr_deref_2835_load_0_req_1 : boolean;
  signal type_cast_2825_inst_ack_0 : boolean;
  signal ptr_deref_2770_load_0_req_0 : boolean;
  signal type_cast_2825_inst_req_0 : boolean;
  signal ptr_deref_2770_load_0_ack_0 : boolean;
  signal ptr_deref_2770_load_0_req_1 : boolean;
  signal ptr_deref_2770_load_0_ack_1 : boolean;
  signal ptr_deref_2851_load_0_ack_1 : boolean;
  signal type_cast_2780_inst_req_0 : boolean;
  signal type_cast_2780_inst_ack_0 : boolean;
  signal type_cast_2780_inst_req_1 : boolean;
  signal type_cast_2780_inst_ack_1 : boolean;
  signal type_cast_3022_inst_req_1 : boolean;
  signal ptr_deref_2835_load_0_ack_0 : boolean;
  signal ptr_deref_2818_load_0_ack_1 : boolean;
  signal ptr_deref_2818_load_0_req_1 : boolean;
  signal ptr_deref_2792_load_0_req_0 : boolean;
  signal ptr_deref_2792_load_0_ack_0 : boolean;
  signal ptr_deref_2792_load_0_req_1 : boolean;
  signal ptr_deref_2792_load_0_ack_1 : boolean;
  signal ptr_deref_2835_load_0_req_0 : boolean;
  signal ptr_deref_2851_load_0_req_1 : boolean;
  signal ptr_deref_2802_load_0_req_0 : boolean;
  signal ptr_deref_2802_load_0_ack_0 : boolean;
  signal ptr_deref_2802_load_0_req_1 : boolean;
  signal ptr_deref_2802_load_0_ack_1 : boolean;
  signal type_cast_3022_inst_ack_1 : boolean;
  signal type_cast_3052_inst_req_0 : boolean;
  signal type_cast_3052_inst_ack_0 : boolean;
  signal type_cast_3052_inst_req_1 : boolean;
  signal type_cast_3052_inst_ack_1 : boolean;
  signal array_obj_ref_3058_index_offset_req_0 : boolean;
  signal array_obj_ref_3058_index_offset_ack_0 : boolean;
  signal array_obj_ref_3058_index_offset_req_1 : boolean;
  signal array_obj_ref_3058_index_offset_ack_1 : boolean;
  signal addr_of_3059_final_reg_req_0 : boolean;
  signal addr_of_3059_final_reg_ack_0 : boolean;
  signal addr_of_3059_final_reg_req_1 : boolean;
  signal addr_of_3059_final_reg_ack_1 : boolean;
  signal ptr_deref_3063_load_0_req_0 : boolean;
  signal ptr_deref_3063_load_0_ack_0 : boolean;
  signal ptr_deref_3063_load_0_req_1 : boolean;
  signal ptr_deref_3063_load_0_ack_1 : boolean;
  signal type_cast_3083_inst_req_0 : boolean;
  signal type_cast_3083_inst_ack_0 : boolean;
  signal type_cast_3083_inst_req_1 : boolean;
  signal type_cast_3083_inst_ack_1 : boolean;
  signal array_obj_ref_3089_index_offset_req_0 : boolean;
  signal array_obj_ref_3089_index_offset_ack_0 : boolean;
  signal array_obj_ref_3089_index_offset_req_1 : boolean;
  signal array_obj_ref_3089_index_offset_ack_1 : boolean;
  signal addr_of_3090_final_reg_req_0 : boolean;
  signal addr_of_3090_final_reg_ack_0 : boolean;
  signal addr_of_3090_final_reg_req_1 : boolean;
  signal addr_of_3090_final_reg_ack_1 : boolean;
  signal ptr_deref_3093_store_0_req_0 : boolean;
  signal ptr_deref_3093_store_0_ack_0 : boolean;
  signal ptr_deref_3093_store_0_req_1 : boolean;
  signal ptr_deref_3093_store_0_ack_1 : boolean;
  signal type_cast_3099_inst_req_0 : boolean;
  signal type_cast_3099_inst_ack_0 : boolean;
  signal type_cast_3099_inst_req_1 : boolean;
  signal type_cast_3099_inst_ack_1 : boolean;
  signal if_stmt_3112_branch_req_0 : boolean;
  signal if_stmt_3112_branch_ack_1 : boolean;
  signal if_stmt_3112_branch_ack_0 : boolean;
  signal type_cast_3136_inst_req_0 : boolean;
  signal type_cast_3136_inst_ack_0 : boolean;
  signal type_cast_3136_inst_req_1 : boolean;
  signal type_cast_3136_inst_ack_1 : boolean;
  signal if_stmt_3143_branch_req_0 : boolean;
  signal if_stmt_3143_branch_ack_1 : boolean;
  signal if_stmt_3143_branch_ack_0 : boolean;
  signal type_cast_3164_inst_req_0 : boolean;
  signal type_cast_3164_inst_ack_0 : boolean;
  signal type_cast_3164_inst_req_1 : boolean;
  signal type_cast_3164_inst_ack_1 : boolean;
  signal type_cast_3184_inst_req_0 : boolean;
  signal type_cast_3184_inst_ack_0 : boolean;
  signal type_cast_3184_inst_req_1 : boolean;
  signal type_cast_3184_inst_ack_1 : boolean;
  signal if_stmt_3191_branch_req_0 : boolean;
  signal if_stmt_3191_branch_ack_1 : boolean;
  signal if_stmt_3191_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_3199_inst_req_0 : boolean;
  signal WPIPE_Block3_done_3199_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_3199_inst_req_1 : boolean;
  signal WPIPE_Block3_done_3199_inst_ack_1 : boolean;
  signal type_cast_2882_inst_req_0 : boolean;
  signal type_cast_2882_inst_ack_0 : boolean;
  signal type_cast_2882_inst_req_1 : boolean;
  signal type_cast_2882_inst_ack_1 : boolean;
  signal phi_stmt_2879_req_0 : boolean;
  signal type_cast_2888_inst_req_0 : boolean;
  signal type_cast_2888_inst_ack_0 : boolean;
  signal type_cast_2888_inst_req_1 : boolean;
  signal type_cast_2888_inst_ack_1 : boolean;
  signal phi_stmt_2885_req_0 : boolean;
  signal type_cast_2884_inst_req_0 : boolean;
  signal type_cast_2884_inst_ack_0 : boolean;
  signal type_cast_2884_inst_req_1 : boolean;
  signal type_cast_2884_inst_ack_1 : boolean;
  signal phi_stmt_2879_req_1 : boolean;
  signal type_cast_2890_inst_req_0 : boolean;
  signal type_cast_2890_inst_ack_0 : boolean;
  signal type_cast_2890_inst_req_1 : boolean;
  signal type_cast_2890_inst_ack_1 : boolean;
  signal phi_stmt_2885_req_1 : boolean;
  signal phi_stmt_2879_ack_0 : boolean;
  signal phi_stmt_2885_ack_0 : boolean;
  signal type_cast_3012_inst_req_0 : boolean;
  signal type_cast_3012_inst_ack_0 : boolean;
  signal type_cast_3012_inst_req_1 : boolean;
  signal type_cast_3012_inst_ack_1 : boolean;
  signal phi_stmt_3006_req_1 : boolean;
  signal phi_stmt_3006_req_0 : boolean;
  signal phi_stmt_3006_ack_0 : boolean;
  signal type_cast_3173_inst_req_0 : boolean;
  signal type_cast_3173_inst_ack_0 : boolean;
  signal type_cast_3173_inst_req_1 : boolean;
  signal type_cast_3173_inst_ack_1 : boolean;
  signal phi_stmt_3168_req_1 : boolean;
  signal type_cast_3179_inst_req_0 : boolean;
  signal type_cast_3179_inst_ack_0 : boolean;
  signal type_cast_3179_inst_req_1 : boolean;
  signal type_cast_3179_inst_ack_1 : boolean;
  signal phi_stmt_3174_req_1 : boolean;
  signal type_cast_3171_inst_req_0 : boolean;
  signal type_cast_3171_inst_ack_0 : boolean;
  signal type_cast_3171_inst_req_1 : boolean;
  signal type_cast_3171_inst_ack_1 : boolean;
  signal phi_stmt_3168_req_0 : boolean;
  signal type_cast_3177_inst_req_0 : boolean;
  signal type_cast_3177_inst_ack_0 : boolean;
  signal type_cast_3177_inst_req_1 : boolean;
  signal type_cast_3177_inst_ack_1 : boolean;
  signal phi_stmt_3174_req_0 : boolean;
  signal phi_stmt_3168_ack_0 : boolean;
  signal phi_stmt_3174_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_7664_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7664_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_7664_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7664_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_7664: Block -- control-path 
    signal convTransposeD_CP_7664_elements: BooleanArray(116 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_7664_elements(0) <= convTransposeD_CP_7664_start;
    convTransposeD_CP_7664_symbol <= convTransposeD_CP_7664_elements(74);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2733/branch_block_stmt_2733__entry__
      -- CP-element group 0: 	 branch_block_stmt_2733/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2733/assign_stmt_2736__entry__
      -- CP-element group 0: 	 branch_block_stmt_2733/assign_stmt_2736/$entry
      -- CP-element group 0: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_Sample/rr
      -- 
    rr_7722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(0), ack => RPIPE_Block3_start_2735_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_Update/cr
      -- 
    ra_7723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2735_inst_ack_0, ack => convTransposeD_CP_7664_elements(1)); -- 
    cr_7727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(1), ack => RPIPE_Block3_start_2735_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	31 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	32 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2:  members (268) 
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876__entry__
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2736__exit__
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2736/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2736/RPIPE_Block3_start_2735_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/word_access_complete/word_0/cr
      -- 
    ca_7728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2735_inst_ack_1, ack => convTransposeD_CP_7664_elements(2)); -- 
    cr_8133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => type_cast_2839_inst_req_1); -- 
    rr_8267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2875_load_0_req_0); -- 
    cr_7972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => type_cast_2806_inst_req_1); -- 
    rr_8039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => LOAD_padding_2821_load_0_req_0); -- 
    cr_8278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2875_load_0_req_1); -- 
    rr_8217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2863_load_0_req_0); -- 
    cr_8050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => LOAD_padding_2821_load_0_req_1); -- 
    cr_8228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2863_load_0_req_1); -- 
    rr_8006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2818_load_0_req_0); -- 
    rr_8167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2851_load_0_req_0); -- 
    rr_7764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2748_load_0_req_0); -- 
    cr_7775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2748_load_0_req_1); -- 
    cr_8069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => type_cast_2825_inst_req_1); -- 
    cr_7794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => type_cast_2758_inst_req_1); -- 
    cr_8114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2835_load_0_req_1); -- 
    rr_7828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2770_load_0_req_0); -- 
    cr_7839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2770_load_0_req_1); -- 
    cr_7858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => type_cast_2780_inst_req_1); -- 
    cr_8017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2818_load_0_req_1); -- 
    rr_7892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2792_load_0_req_0); -- 
    cr_7903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2792_load_0_req_1); -- 
    rr_8103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2835_load_0_req_0); -- 
    cr_8178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2851_load_0_req_1); -- 
    rr_7942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2802_load_0_req_0); -- 
    cr_7953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2802_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Sample/word_access_start/word_0/ra
      -- 
    ra_7765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2748_load_0_ack_0, ack => convTransposeD_CP_7664_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/ptr_deref_2748_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/ptr_deref_2748_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/ptr_deref_2748_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2748_Update/ptr_deref_2748_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_Sample/rr
      -- 
    ca_7776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2748_load_0_ack_1, ack => convTransposeD_CP_7664_elements(4)); -- 
    rr_7789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(4), ack => type_cast_2758_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_Sample/ra
      -- 
    ra_7790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2758_inst_ack_0, ack => convTransposeD_CP_7664_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	33 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2758_Update/ca
      -- 
    ca_7795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2758_inst_ack_1, ack => convTransposeD_CP_7664_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Sample/word_access_start/word_0/ra
      -- 
    ra_7829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2770_load_0_ack_0, ack => convTransposeD_CP_7664_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/ptr_deref_2770_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/ptr_deref_2770_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/ptr_deref_2770_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2770_Update/ptr_deref_2770_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_Sample/rr
      -- 
    ca_7840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2770_load_0_ack_1, ack => convTransposeD_CP_7664_elements(8)); -- 
    rr_7853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(8), ack => type_cast_2780_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_Sample/ra
      -- 
    ra_7854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2780_inst_ack_0, ack => convTransposeD_CP_7664_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	33 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2780_Update/ca
      -- 
    ca_7859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2780_inst_ack_1, ack => convTransposeD_CP_7664_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Sample/word_access_start/word_0/ra
      -- 
    ra_7893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2792_load_0_ack_0, ack => convTransposeD_CP_7664_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	33 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/ptr_deref_2792_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/ptr_deref_2792_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/ptr_deref_2792_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2792_Update/ptr_deref_2792_Merge/merge_ack
      -- 
    ca_7904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2792_load_0_ack_1, ack => convTransposeD_CP_7664_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Sample/word_access_start/word_0/ra
      -- 
    ra_7943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2802_load_0_ack_0, ack => convTransposeD_CP_7664_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/ptr_deref_2802_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/ptr_deref_2802_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/ptr_deref_2802_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2802_Update/ptr_deref_2802_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_sample_start_
      -- 
    ca_7954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2802_load_0_ack_1, ack => convTransposeD_CP_7664_elements(14)); -- 
    rr_7967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(14), ack => type_cast_2806_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_sample_completed_
      -- 
    ra_7968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2806_inst_ack_0, ack => convTransposeD_CP_7664_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	33 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2806_update_completed_
      -- 
    ca_7973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2806_inst_ack_1, ack => convTransposeD_CP_7664_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Sample/word_access_start/word_0/ra
      -- CP-element group 17: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Sample/word_access_start/word_0/$exit
      -- 
    ra_8007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2818_load_0_ack_0, ack => convTransposeD_CP_7664_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	33 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/ptr_deref_2818_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/ptr_deref_2818_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/ptr_deref_2818_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/ptr_deref_2818_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2818_Update/word_access_complete/word_0/$exit
      -- 
    ca_8018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2818_load_0_ack_1, ack => convTransposeD_CP_7664_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Sample/word_access_start/word_0/ra
      -- CP-element group 19: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_sample_completed_
      -- 
    ra_8040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2821_load_0_ack_0, ack => convTransposeD_CP_7664_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/LOAD_padding_2821_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/LOAD_padding_2821_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/LOAD_padding_2821_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/LOAD_padding_2821_Update/LOAD_padding_2821_Merge/$entry
      -- 
    ca_8051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2821_load_0_ack_1, ack => convTransposeD_CP_7664_elements(20)); -- 
    rr_8064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(20), ack => type_cast_2825_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_sample_completed_
      -- 
    ra_8065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2825_inst_ack_0, ack => convTransposeD_CP_7664_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	33 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2825_update_completed_
      -- 
    ca_8070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2825_inst_ack_1, ack => convTransposeD_CP_7664_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Sample/word_access_start/word_0/ra
      -- CP-element group 23: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Sample/word_access_start/word_0/$exit
      -- 
    ra_8104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2835_load_0_ack_0, ack => convTransposeD_CP_7664_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (12) 
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/ptr_deref_2835_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/ptr_deref_2835_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/ptr_deref_2835_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/ptr_deref_2835_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2835_Update/$exit
      -- 
    ca_8115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2835_load_0_ack_1, ack => convTransposeD_CP_7664_elements(24)); -- 
    rr_8128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(24), ack => type_cast_2839_inst_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_sample_completed_
      -- 
    ra_8129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2839_inst_ack_0, ack => convTransposeD_CP_7664_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	33 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/type_cast_2839_update_completed_
      -- 
    ca_8134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2839_inst_ack_1, ack => convTransposeD_CP_7664_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Sample/word_access_start/word_0/ra
      -- CP-element group 27: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_sample_completed_
      -- 
    ra_8168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2851_load_0_ack_0, ack => convTransposeD_CP_7664_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	33 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/ptr_deref_2851_Merge/merge_ack
      -- CP-element group 28: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/ptr_deref_2851_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/ptr_deref_2851_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/ptr_deref_2851_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2851_update_completed_
      -- 
    ca_8179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2851_load_0_ack_1, ack => convTransposeD_CP_7664_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Sample/word_access_start/word_0/ra
      -- 
    ra_8218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2863_load_0_ack_0, ack => convTransposeD_CP_7664_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/ptr_deref_2863_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/ptr_deref_2863_Merge/merge_ack
      -- CP-element group 30: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/ptr_deref_2863_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/ptr_deref_2863_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2863_Update/$exit
      -- 
    ca_8229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2863_load_0_ack_1, ack => convTransposeD_CP_7664_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	2 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Sample/word_access_start/word_0/ra
      -- CP-element group 31: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Sample/word_access_start/$exit
      -- 
    ra_8268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2875_load_0_ack_0, ack => convTransposeD_CP_7664_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	2 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/word_access_complete/$exit
      -- CP-element group 32: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/ptr_deref_2875_Merge/$entry
      -- CP-element group 32: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/ptr_deref_2875_Merge/$exit
      -- CP-element group 32: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/ptr_deref_2875_Merge/merge_ack
      -- CP-element group 32: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/word_access_complete/word_0/ca
      -- CP-element group 32: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/ptr_deref_2875_Update/ptr_deref_2875_Merge/merge_req
      -- 
    ca_8279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2875_load_0_ack_1, ack => convTransposeD_CP_7664_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  place  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	22 
    -- CP-element group 33: 	28 
    -- CP-element group 33: 	18 
    -- CP-element group 33: 	32 
    -- CP-element group 33: 	26 
    -- CP-element group 33: 	30 
    -- CP-element group 33: 	6 
    -- CP-element group 33: 	10 
    -- CP-element group 33: 	12 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	75 
    -- CP-element group 33: 	76 
    -- CP-element group 33: 	78 
    -- CP-element group 33: 	79 
    -- CP-element group 33:  members (20) 
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter
      -- CP-element group 33: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876__exit__
      -- CP-element group 33: 	 branch_block_stmt_2733/assign_stmt_2745_to_assign_stmt_2876/$exit
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/SplitProtocol/Update/cr
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Update/cr
      -- 
    rr_8713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(33), ack => type_cast_2882_inst_req_0); -- 
    cr_8718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(33), ack => type_cast_2882_inst_req_1); -- 
    rr_8736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(33), ack => type_cast_2888_inst_req_0); -- 
    cr_8741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(33), ack => type_cast_2888_inst_req_1); -- 
    convTransposeD_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(16) & convTransposeD_CP_7664_elements(22) & convTransposeD_CP_7664_elements(28) & convTransposeD_CP_7664_elements(18) & convTransposeD_CP_7664_elements(32) & convTransposeD_CP_7664_elements(26) & convTransposeD_CP_7664_elements(30) & convTransposeD_CP_7664_elements(6) & convTransposeD_CP_7664_elements(10) & convTransposeD_CP_7664_elements(12);
      gj_convTransposeD_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	92 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_Sample/ra
      -- 
    ra_8296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2895_inst_ack_0, ack => convTransposeD_CP_7664_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	92 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_Update/$exit
      -- 
    ca_8301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2895_inst_ack_1, ack => convTransposeD_CP_7664_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	92 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_Sample/ra
      -- 
    ra_8310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2900_inst_ack_0, ack => convTransposeD_CP_7664_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_Update/ca
      -- 
    ca_8315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2900_inst_ack_1, ack => convTransposeD_CP_7664_elements(37)); -- 
    -- CP-element group 38:  join  transition  place  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	96 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/$exit
      -- CP-element group 38: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003__exit__
      -- CP-element group 38: 	 branch_block_stmt_2733/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 38: 	 branch_block_stmt_2733/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_2733/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3006/$entry
      -- CP-element group 38: 	 branch_block_stmt_2733/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/$entry
      -- 
    convTransposeD_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(37) & convTransposeD_CP_7664_elements(35);
      gj_convTransposeD_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	98 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_Sample/ra
      -- 
    ra_8327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3022_inst_ack_0, ack => convTransposeD_CP_7664_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	98 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	49 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_Sample/rr
      -- CP-element group 40: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_Sample/rr
      -- 
    ca_8332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3022_inst_ack_1, ack => convTransposeD_CP_7664_elements(40)); -- 
    rr_8450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(40), ack => type_cast_3083_inst_req_0); -- 
    rr_8340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(40), ack => type_cast_3052_inst_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_Sample/ra
      -- 
    ra_8341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3052_inst_ack_0, ack => convTransposeD_CP_7664_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	98 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (16) 
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_resized_1
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_scaled_1
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_computed_1
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_resize_1/$entry
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_resize_1/$exit
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_resize_1/index_resize_req
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_resize_1/index_resize_ack
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_scale_1/$entry
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_scale_1/$exit
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_scale_1/scale_rename_req
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_index_scale_1/scale_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_final_index_sum_regn_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_final_index_sum_regn_Sample/req
      -- 
    ca_8346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3052_inst_ack_1, ack => convTransposeD_CP_7664_elements(42)); -- 
    req_8371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(42), ack => array_obj_ref_3058_index_offset_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	60 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_final_index_sum_regn_sample_complete
      -- CP-element group 43: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_final_index_sum_regn_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_final_index_sum_regn_Sample/ack
      -- 
    ack_8372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3058_index_offset_ack_0, ack => convTransposeD_CP_7664_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	98 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (11) 
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_offset_calculated
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_final_index_sum_regn_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_final_index_sum_regn_Update/ack
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_request/$entry
      -- CP-element group 44: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_request/req
      -- 
    ack_8377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3058_index_offset_ack_1, ack => convTransposeD_CP_7664_elements(44)); -- 
    req_8386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(44), ack => addr_of_3059_final_reg_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_request/$exit
      -- CP-element group 45: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_request/ack
      -- 
    ack_8387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3059_final_reg_ack_0, ack => convTransposeD_CP_7664_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	98 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (24) 
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_complete/ack
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_base_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_word_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_root_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_base_address_resized
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_base_addr_resize/$entry
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_base_addr_resize/$exit
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_base_addr_resize/base_resize_req
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_base_addr_resize/base_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_base_plus_offset/$entry
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_base_plus_offset/$exit
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_base_plus_offset/sum_rename_req
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_base_plus_offset/sum_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_word_addrgen/$entry
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_word_addrgen/$exit
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_word_addrgen/root_register_req
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_word_addrgen/root_register_ack
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Sample/word_access_start/$entry
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Sample/word_access_start/word_0/$entry
      -- CP-element group 46: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Sample/word_access_start/word_0/rr
      -- 
    ack_8392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3059_final_reg_ack_1, ack => convTransposeD_CP_7664_elements(46)); -- 
    rr_8425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(46), ack => ptr_deref_3063_load_0_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Sample/word_access_start/$exit
      -- CP-element group 47: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Sample/word_access_start/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Sample/word_access_start/word_0/ra
      -- 
    ra_8426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3063_load_0_ack_0, ack => convTransposeD_CP_7664_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	98 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	55 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/word_access_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/word_access_complete/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/word_access_complete/word_0/ca
      -- CP-element group 48: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/ptr_deref_3063_Merge/$entry
      -- CP-element group 48: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/ptr_deref_3063_Merge/$exit
      -- CP-element group 48: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/ptr_deref_3063_Merge/merge_req
      -- CP-element group 48: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/ptr_deref_3063_Merge/merge_ack
      -- 
    ca_8437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3063_load_0_ack_1, ack => convTransposeD_CP_7664_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	40 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_Sample/ra
      -- 
    ra_8451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3083_inst_ack_0, ack => convTransposeD_CP_7664_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	98 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (16) 
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_resized_1
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_scaled_1
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_computed_1
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_resize_1/$entry
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_resize_1/$exit
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_resize_1/index_resize_req
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_resize_1/index_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_scale_1/$entry
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_scale_1/$exit
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_scale_1/scale_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_index_scale_1/scale_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_final_index_sum_regn_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_final_index_sum_regn_Sample/req
      -- 
    ca_8456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3083_inst_ack_1, ack => convTransposeD_CP_7664_elements(50)); -- 
    req_8481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(50), ack => array_obj_ref_3089_index_offset_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	60 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_final_index_sum_regn_sample_complete
      -- CP-element group 51: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_final_index_sum_regn_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_final_index_sum_regn_Sample/ack
      -- 
    ack_8482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3089_index_offset_ack_0, ack => convTransposeD_CP_7664_elements(51)); -- 
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	98 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (11) 
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_request/$entry
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_offset_calculated
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_final_index_sum_regn_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_final_index_sum_regn_Update/ack
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_request/req
      -- 
    ack_8487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3089_index_offset_ack_1, ack => convTransposeD_CP_7664_elements(52)); -- 
    req_8496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(52), ack => addr_of_3090_final_reg_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_request/$exit
      -- CP-element group 53: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_request/ack
      -- 
    ack_8497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3090_final_reg_ack_0, ack => convTransposeD_CP_7664_elements(53)); -- 
    -- CP-element group 54:  fork  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	98 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (19) 
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_complete/$exit
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_complete/ack
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_base_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_word_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_root_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_base_address_resized
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_base_addr_resize/$entry
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_base_addr_resize/$exit
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_base_addr_resize/base_resize_req
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_base_addr_resize/base_resize_ack
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_base_plus_offset/$entry
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_base_plus_offset/$exit
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_base_plus_offset/sum_rename_req
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_base_plus_offset/sum_rename_ack
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_word_addrgen/$entry
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_word_addrgen/$exit
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_word_addrgen/root_register_req
      -- CP-element group 54: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_word_addrgen/root_register_ack
      -- 
    ack_8502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3090_final_reg_ack_1, ack => convTransposeD_CP_7664_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	48 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/ptr_deref_3093_Split/$entry
      -- CP-element group 55: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/ptr_deref_3093_Split/$exit
      -- CP-element group 55: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/ptr_deref_3093_Split/split_req
      -- CP-element group 55: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/ptr_deref_3093_Split/split_ack
      -- CP-element group 55: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/word_access_start/word_0/rr
      -- 
    rr_8540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(55), ack => ptr_deref_3093_store_0_req_0); -- 
    convTransposeD_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(54) & convTransposeD_CP_7664_elements(48);
      gj_convTransposeD_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Sample/word_access_start/word_0/ra
      -- 
    ra_8541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3093_store_0_ack_0, ack => convTransposeD_CP_7664_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	98 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	60 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Update/word_access_complete/word_0/ca
      -- 
    ca_8552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3093_store_0_ack_1, ack => convTransposeD_CP_7664_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	98 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_Sample/ra
      -- 
    ra_8561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3099_inst_ack_0, ack => convTransposeD_CP_7664_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	98 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_Update/ca
      -- 
    ca_8566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3099_inst_ack_1, ack => convTransposeD_CP_7664_elements(59)); -- 
    -- CP-element group 60:  branch  join  transition  place  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	57 
    -- CP-element group 60: 	43 
    -- CP-element group 60: 	59 
    -- CP-element group 60: 	51 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (10) 
      -- CP-element group 60: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/$exit
      -- CP-element group 60: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111__exit__
      -- CP-element group 60: 	 branch_block_stmt_2733/if_stmt_3112__entry__
      -- CP-element group 60: 	 branch_block_stmt_2733/R_cmp_3113_place
      -- CP-element group 60: 	 branch_block_stmt_2733/if_stmt_3112_dead_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_2733/if_stmt_3112_eval_test/$entry
      -- CP-element group 60: 	 branch_block_stmt_2733/if_stmt_3112_eval_test/$exit
      -- CP-element group 60: 	 branch_block_stmt_2733/if_stmt_3112_eval_test/branch_req
      -- CP-element group 60: 	 branch_block_stmt_2733/if_stmt_3112_if_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_2733/if_stmt_3112_else_link/$entry
      -- 
    branch_req_8574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(60), ack => if_stmt_3112_branch_req_0); -- 
    convTransposeD_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(57) & convTransposeD_CP_7664_elements(43) & convTransposeD_CP_7664_elements(59) & convTransposeD_CP_7664_elements(51);
      gj_convTransposeD_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	93 
    -- CP-element group 61: 	94 
    -- CP-element group 61:  members (24) 
      -- CP-element group 61: 	 branch_block_stmt_2733/whilex_xbody_ifx_xthen
      -- CP-element group 61: 	 branch_block_stmt_2733/merge_stmt_3118__exit__
      -- CP-element group 61: 	 branch_block_stmt_2733/assign_stmt_3124__entry__
      -- CP-element group 61: 	 branch_block_stmt_2733/assign_stmt_3124__exit__
      -- CP-element group 61: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody
      -- CP-element group 61: 	 branch_block_stmt_2733/if_stmt_3112_if_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_2733/if_stmt_3112_if_link/if_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_2733/assign_stmt_3124/$entry
      -- CP-element group 61: 	 branch_block_stmt_2733/assign_stmt_3124/$exit
      -- CP-element group 61: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/$entry
      -- CP-element group 61: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/$entry
      -- CP-element group 61: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/SplitProtocol/Update/cr
      -- CP-element group 61: 	 branch_block_stmt_2733/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2733/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_2733/merge_stmt_3118_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_2733/merge_stmt_3118_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_2733/merge_stmt_3118_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_2733/merge_stmt_3118_PhiAck/dummy
      -- 
    if_choice_transition_8579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3112_branch_ack_1, ack => convTransposeD_CP_7664_elements(61)); -- 
    rr_8817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(61), ack => type_cast_3012_inst_req_0); -- 
    cr_8822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(61), ack => type_cast_3012_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (18) 
      -- CP-element group 62: 	 branch_block_stmt_2733/whilex_xbody_ifx_xelse
      -- CP-element group 62: 	 branch_block_stmt_2733/merge_stmt_3126__exit__
      -- CP-element group 62: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142__entry__
      -- CP-element group 62: 	 branch_block_stmt_2733/if_stmt_3112_else_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_2733/if_stmt_3112_else_link/else_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/$entry
      -- CP-element group 62: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_2733/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_2733/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_2733/merge_stmt_3126_PhiReqMerge
      -- CP-element group 62: 	 branch_block_stmt_2733/merge_stmt_3126_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_2733/merge_stmt_3126_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_2733/merge_stmt_3126_PhiAck/dummy
      -- 
    else_choice_transition_8583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3112_branch_ack_0, ack => convTransposeD_CP_7664_elements(62)); -- 
    rr_8599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(62), ack => type_cast_3136_inst_req_0); -- 
    cr_8604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(62), ack => type_cast_3136_inst_req_1); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_Sample/ra
      -- 
    ra_8600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3136_inst_ack_0, ack => convTransposeD_CP_7664_elements(63)); -- 
    -- CP-element group 64:  branch  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142__exit__
      -- CP-element group 64: 	 branch_block_stmt_2733/if_stmt_3143__entry__
      -- CP-element group 64: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/$exit
      -- CP-element group 64: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2733/assign_stmt_3132_to_assign_stmt_3142/type_cast_3136_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2733/if_stmt_3143_dead_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_2733/if_stmt_3143_eval_test/$entry
      -- CP-element group 64: 	 branch_block_stmt_2733/if_stmt_3143_eval_test/$exit
      -- CP-element group 64: 	 branch_block_stmt_2733/if_stmt_3143_eval_test/branch_req
      -- CP-element group 64: 	 branch_block_stmt_2733/R_cmp81_3144_place
      -- CP-element group 64: 	 branch_block_stmt_2733/if_stmt_3143_if_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_2733/if_stmt_3143_else_link/$entry
      -- 
    ca_8605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3136_inst_ack_1, ack => convTransposeD_CP_7664_elements(64)); -- 
    branch_req_8613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(64), ack => if_stmt_3143_branch_req_0); -- 
    -- CP-element group 65:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (18) 
      -- CP-element group 65: 	 branch_block_stmt_2733/merge_stmt_3149__exit__
      -- CP-element group 65: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165__entry__
      -- CP-element group 65: 	 branch_block_stmt_2733/if_stmt_3143_if_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_2733/if_stmt_3143_if_link/if_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_2733/ifx_xelse_ifx_xthen83
      -- CP-element group 65: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/$entry
      -- CP-element group 65: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_update_start_
      -- CP-element group 65: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_2733/ifx_xelse_ifx_xthen83_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_2733/ifx_xelse_ifx_xthen83_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_2733/merge_stmt_3149_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_2733/merge_stmt_3149_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_2733/merge_stmt_3149_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_2733/merge_stmt_3149_PhiAck/dummy
      -- 
    if_choice_transition_8618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3143_branch_ack_1, ack => convTransposeD_CP_7664_elements(65)); -- 
    rr_8635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(65), ack => type_cast_3164_inst_req_0); -- 
    cr_8640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(65), ack => type_cast_3164_inst_req_1); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	99 
    -- CP-element group 66: 	100 
    -- CP-element group 66: 	102 
    -- CP-element group 66: 	103 
    -- CP-element group 66:  members (20) 
      -- CP-element group 66: 	 branch_block_stmt_2733/if_stmt_3143_else_link/$exit
      -- CP-element group 66: 	 branch_block_stmt_2733/if_stmt_3143_else_link/else_choice_transition
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3143_branch_ack_0, ack => convTransposeD_CP_7664_elements(66)); -- 
    rr_8891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(66), ack => type_cast_3173_inst_req_0); -- 
    cr_8896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(66), ack => type_cast_3173_inst_req_1); -- 
    rr_8914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(66), ack => type_cast_3179_inst_req_0); -- 
    cr_8919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(66), ack => type_cast_3179_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_Sample/ra
      -- 
    ra_8636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3164_inst_ack_0, ack => convTransposeD_CP_7664_elements(67)); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	106 
    -- CP-element group 68: 	107 
    -- CP-element group 68: 	109 
    -- CP-element group 68: 	110 
    -- CP-element group 68:  members (23) 
      -- CP-element group 68: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165__exit__
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend
      -- CP-element group 68: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/$exit
      -- CP-element group 68: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2733/assign_stmt_3155_to_assign_stmt_3165/type_cast_3164_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/SplitProtocol/Update/cr
      -- 
    ca_8641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3164_inst_ack_1, ack => convTransposeD_CP_7664_elements(68)); -- 
    rr_8940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(68), ack => type_cast_3171_inst_req_0); -- 
    cr_8945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(68), ack => type_cast_3171_inst_req_1); -- 
    rr_8963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(68), ack => type_cast_3177_inst_req_0); -- 
    cr_8968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(68), ack => type_cast_3177_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	116 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_Sample/ra
      -- 
    ra_8653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3184_inst_ack_0, ack => convTransposeD_CP_7664_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	116 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190__exit__
      -- CP-element group 70: 	 branch_block_stmt_2733/if_stmt_3191__entry__
      -- CP-element group 70: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/$exit
      -- CP-element group 70: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2733/if_stmt_3191_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2733/if_stmt_3191_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2733/if_stmt_3191_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2733/if_stmt_3191_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2733/R_cmp92_3192_place
      -- CP-element group 70: 	 branch_block_stmt_2733/if_stmt_3191_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2733/if_stmt_3191_else_link/$entry
      -- 
    ca_8658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3184_inst_ack_1, ack => convTransposeD_CP_7664_elements(70)); -- 
    branch_req_8666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(70), ack => if_stmt_3191_branch_req_0); -- 
    -- CP-element group 71:  merge  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2733/merge_stmt_3197__exit__
      -- CP-element group 71: 	 branch_block_stmt_2733/assign_stmt_3201__entry__
      -- CP-element group 71: 	 branch_block_stmt_2733/if_stmt_3191_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2733/if_stmt_3191_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2733/ifx_xend_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2733/assign_stmt_3201/$entry
      -- CP-element group 71: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2733/ifx_xend_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2733/ifx_xend_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2733/merge_stmt_3197_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2733/merge_stmt_3197_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2733/merge_stmt_3197_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2733/merge_stmt_3197_PhiAck/dummy
      -- 
    if_choice_transition_8671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3191_branch_ack_1, ack => convTransposeD_CP_7664_elements(71)); -- 
    req_8688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(71), ack => WPIPE_Block3_done_3199_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	82 
    -- CP-element group 72: 	83 
    -- CP-element group 72: 	85 
    -- CP-element group 72: 	86 
    -- CP-element group 72:  members (20) 
      -- CP-element group 72: 	 branch_block_stmt_2733/if_stmt_3191_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2733/if_stmt_3191_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3191_branch_ack_0, ack => convTransposeD_CP_7664_elements(72)); -- 
    rr_8762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(72), ack => type_cast_2884_inst_req_0); -- 
    cr_8767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(72), ack => type_cast_2884_inst_req_1); -- 
    rr_8785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(72), ack => type_cast_2890_inst_req_0); -- 
    cr_8790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(72), ack => type_cast_2890_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_Update/req
      -- 
    ack_8689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3199_inst_ack_0, ack => convTransposeD_CP_7664_elements(73)); -- 
    req_8693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(73), ack => WPIPE_Block3_done_3199_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 branch_block_stmt_2733/branch_block_stmt_2733__exit__
      -- CP-element group 74: 	 branch_block_stmt_2733/$exit
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2733/assign_stmt_3201__exit__
      -- CP-element group 74: 	 branch_block_stmt_2733/return__
      -- CP-element group 74: 	 branch_block_stmt_2733/merge_stmt_3203__exit__
      -- CP-element group 74: 	 branch_block_stmt_2733/assign_stmt_3201/$exit
      -- CP-element group 74: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2733/assign_stmt_3201/WPIPE_Block3_done_3199_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2733/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2733/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2733/merge_stmt_3203_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2733/merge_stmt_3203_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2733/merge_stmt_3203_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2733/merge_stmt_3203_PhiAck/dummy
      -- 
    ack_8694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3199_inst_ack_1, ack => convTransposeD_CP_7664_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	33 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/SplitProtocol/Sample/ra
      -- 
    ra_8714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2882_inst_ack_0, ack => convTransposeD_CP_7664_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	33 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/SplitProtocol/Update/ca
      -- 
    ca_8719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2882_inst_ack_1, ack => convTransposeD_CP_7664_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/$exit
      -- CP-element group 77: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/$exit
      -- CP-element group 77: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2882/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_req
      -- 
    phi_stmt_2879_req_8720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2879_req_8720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(77), ack => phi_stmt_2879_req_0); -- 
    convTransposeD_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(75) & convTransposeD_CP_7664_elements(76);
      gj_convTransposeD_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	33 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Sample/ra
      -- 
    ra_8737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2888_inst_ack_0, ack => convTransposeD_CP_7664_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	33 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/Update/ca
      -- 
    ca_8742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2888_inst_ack_1, ack => convTransposeD_CP_7664_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/$exit
      -- CP-element group 80: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/$exit
      -- CP-element group 80: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2888/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_req
      -- 
    phi_stmt_2885_req_8743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2885_req_8743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(80), ack => phi_stmt_2885_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(78) & convTransposeD_CP_7664_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	89 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2733/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(77) & convTransposeD_CP_7664_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	72 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/SplitProtocol/Sample/ra
      -- 
    ra_8763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2884_inst_ack_0, ack => convTransposeD_CP_7664_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	72 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/SplitProtocol/Update/ca
      -- 
    ca_8768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2884_inst_ack_1, ack => convTransposeD_CP_7664_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	88 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/$exit
      -- CP-element group 84: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/$exit
      -- CP-element group 84: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_sources/type_cast_2884/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2879/phi_stmt_2879_req
      -- 
    phi_stmt_2879_req_8769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2879_req_8769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(84), ack => phi_stmt_2879_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(82) & convTransposeD_CP_7664_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	72 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/SplitProtocol/Sample/ra
      -- 
    ra_8786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2890_inst_ack_0, ack => convTransposeD_CP_7664_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	72 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/SplitProtocol/Update/ca
      -- 
    ca_8791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2890_inst_ack_1, ack => convTransposeD_CP_7664_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/$exit
      -- CP-element group 87: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/$exit
      -- CP-element group 87: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_sources/type_cast_2890/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2885/phi_stmt_2885_req
      -- 
    phi_stmt_2885_req_8792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2885_req_8792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(87), ack => phi_stmt_2885_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(85) & convTransposeD_CP_7664_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	84 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2733/ifx_xend_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(84) & convTransposeD_CP_7664_elements(87);
      gj_convTransposeD_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  merge  fork  transition  place  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	81 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2733/merge_stmt_2878_PhiReqMerge
      -- CP-element group 89: 	 branch_block_stmt_2733/merge_stmt_2878_PhiAck/$entry
      -- 
    convTransposeD_CP_7664_elements(89) <= OrReduce(convTransposeD_CP_7664_elements(81) & convTransposeD_CP_7664_elements(88));
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2733/merge_stmt_2878_PhiAck/phi_stmt_2879_ack
      -- 
    phi_stmt_2879_ack_8797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2879_ack_0, ack => convTransposeD_CP_7664_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_2733/merge_stmt_2878_PhiAck/phi_stmt_2885_ack
      -- 
    phi_stmt_2885_ack_8798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2885_ack_0, ack => convTransposeD_CP_7664_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  place  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	36 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	34 
    -- CP-element group 92: 	35 
    -- CP-element group 92:  members (16) 
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/$entry
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2733/merge_stmt_2878__exit__
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003__entry__
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2895_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2733/assign_stmt_2896_to_assign_stmt_3003/type_cast_2900_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2733/merge_stmt_2878_PhiAck/$exit
      -- 
    rr_8309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(92), ack => type_cast_2900_inst_req_0); -- 
    rr_8295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(92), ack => type_cast_2895_inst_req_0); -- 
    cr_8300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(92), ack => type_cast_2895_inst_req_1); -- 
    cr_8314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(92), ack => type_cast_2900_inst_req_1); -- 
    convTransposeD_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(90) & convTransposeD_CP_7664_elements(91);
      gj_convTransposeD_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	61 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/SplitProtocol/Sample/ra
      -- 
    ra_8818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3012_inst_ack_0, ack => convTransposeD_CP_7664_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	61 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/SplitProtocol/Update/ca
      -- 
    ca_8823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3012_inst_ack_1, ack => convTransposeD_CP_7664_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 95: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/$exit
      -- CP-element group 95: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/$exit
      -- CP-element group 95: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3012/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_2733/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_req
      -- 
    phi_stmt_3006_req_8824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3006_req_8824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(95), ack => phi_stmt_3006_req_1); -- 
    convTransposeD_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(93) & convTransposeD_CP_7664_elements(94);
      gj_convTransposeD_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  transition  output  delay-element  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	38 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_2733/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 96: 	 branch_block_stmt_2733/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3006/$exit
      -- CP-element group 96: 	 branch_block_stmt_2733/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_2733/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_sources/type_cast_3010_konst_delay_trans
      -- CP-element group 96: 	 branch_block_stmt_2733/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3006/phi_stmt_3006_req
      -- 
    phi_stmt_3006_req_8835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3006_req_8835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(96), ack => phi_stmt_3006_req_0); -- 
    -- Element group convTransposeD_CP_7664_elements(96) is a control-delay.
    cp_element_96_delay: control_delay_element  generic map(name => " 96_delay", delay_value => 1)  port map(req => convTransposeD_CP_7664_elements(38), ack => convTransposeD_CP_7664_elements(96), clk => clk, reset =>reset);
    -- CP-element group 97:  merge  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_2733/merge_stmt_3005_PhiReqMerge
      -- CP-element group 97: 	 branch_block_stmt_2733/merge_stmt_3005_PhiAck/$entry
      -- 
    convTransposeD_CP_7664_elements(97) <= OrReduce(convTransposeD_CP_7664_elements(95) & convTransposeD_CP_7664_elements(96));
    -- CP-element group 98:  fork  transition  place  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	57 
    -- CP-element group 98: 	54 
    -- CP-element group 98: 	39 
    -- CP-element group 98: 	50 
    -- CP-element group 98: 	58 
    -- CP-element group 98: 	59 
    -- CP-element group 98: 	52 
    -- CP-element group 98: 	48 
    -- CP-element group 98: 	46 
    -- CP-element group 98: 	40 
    -- CP-element group 98: 	42 
    -- CP-element group 98: 	44 
    -- CP-element group 98:  members (45) 
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_2733/merge_stmt_3005__exit__
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111__entry__
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3022_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3052_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_final_index_sum_regn_update_start
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_final_index_sum_regn_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3058_final_index_sum_regn_Update/req
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3059_complete/req
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/word_access_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/word_access_complete/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3063_Update/word_access_complete/word_0/cr
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3083_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_final_index_sum_regn_update_start
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_final_index_sum_regn_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/array_obj_ref_3089_final_index_sum_regn_Update/req
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/addr_of_3090_complete/req
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Update/word_access_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Update/word_access_complete/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/ptr_deref_3093_Update/word_access_complete/word_0/cr
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2733/assign_stmt_3019_to_assign_stmt_3111/type_cast_3099_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2733/merge_stmt_3005_PhiAck/$exit
      -- CP-element group 98: 	 branch_block_stmt_2733/merge_stmt_3005_PhiAck/phi_stmt_3006_ack
      -- 
    phi_stmt_3006_ack_8840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3006_ack_0, ack => convTransposeD_CP_7664_elements(98)); -- 
    rr_8326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3022_inst_req_0); -- 
    cr_8331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3022_inst_req_1); -- 
    cr_8345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3052_inst_req_1); -- 
    req_8376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => array_obj_ref_3058_index_offset_req_1); -- 
    req_8391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => addr_of_3059_final_reg_req_1); -- 
    cr_8436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => ptr_deref_3063_load_0_req_1); -- 
    cr_8455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3083_inst_req_1); -- 
    req_8486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => array_obj_ref_3089_index_offset_req_1); -- 
    req_8501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => addr_of_3090_final_reg_req_1); -- 
    cr_8551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => ptr_deref_3093_store_0_req_1); -- 
    rr_8560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3099_inst_req_0); -- 
    cr_8565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3099_inst_req_1); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	66 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/SplitProtocol/Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/SplitProtocol/Sample/ra
      -- 
    ra_8892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3173_inst_ack_0, ack => convTransposeD_CP_7664_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	66 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/SplitProtocol/Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/SplitProtocol/Update/ca
      -- 
    ca_8897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3173_inst_ack_1, ack => convTransposeD_CP_7664_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	105 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/$exit
      -- CP-element group 101: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/$exit
      -- CP-element group 101: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3173/SplitProtocol/$exit
      -- CP-element group 101: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_req
      -- 
    phi_stmt_3168_req_8898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3168_req_8898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(101), ack => phi_stmt_3168_req_1); -- 
    convTransposeD_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(99) & convTransposeD_CP_7664_elements(100);
      gj_convTransposeD_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	66 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/SplitProtocol/Sample/ra
      -- 
    ra_8915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3179_inst_ack_0, ack => convTransposeD_CP_7664_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/SplitProtocol/Update/ca
      -- 
    ca_8920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3179_inst_ack_1, ack => convTransposeD_CP_7664_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/$exit
      -- CP-element group 104: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/$exit
      -- CP-element group 104: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3179/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_req
      -- 
    phi_stmt_3174_req_8921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3174_req_8921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(104), ack => phi_stmt_3174_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(102) & convTransposeD_CP_7664_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	101 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	113 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_2733/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(101) & convTransposeD_CP_7664_elements(104);
      gj_convTransposeD_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	68 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/SplitProtocol/Sample/ra
      -- 
    ra_8941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3171_inst_ack_0, ack => convTransposeD_CP_7664_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	68 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/SplitProtocol/Update/ca
      -- 
    ca_8946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3171_inst_ack_1, ack => convTransposeD_CP_7664_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/$exit
      -- CP-element group 108: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/$exit
      -- CP-element group 108: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_sources/type_cast_3171/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3168/phi_stmt_3168_req
      -- 
    phi_stmt_3168_req_8947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3168_req_8947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(108), ack => phi_stmt_3168_req_0); -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(106) & convTransposeD_CP_7664_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	68 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/SplitProtocol/Sample/ra
      -- 
    ra_8964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3177_inst_ack_0, ack => convTransposeD_CP_7664_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	68 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/SplitProtocol/Update/ca
      -- 
    ca_8969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3177_inst_ack_1, ack => convTransposeD_CP_7664_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/$exit
      -- CP-element group 111: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/$exit
      -- CP-element group 111: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_sources/type_cast_3177/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3174/phi_stmt_3174_req
      -- 
    phi_stmt_3174_req_8970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3174_req_8970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(111), ack => phi_stmt_3174_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(109) & convTransposeD_CP_7664_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2733/ifx_xthen83_ifx_xend_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(108) & convTransposeD_CP_7664_elements(111);
      gj_convTransposeD_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  merge  fork  transition  place  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	105 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2733/merge_stmt_3167_PhiReqMerge
      -- CP-element group 113: 	 branch_block_stmt_2733/merge_stmt_3167_PhiAck/$entry
      -- 
    convTransposeD_CP_7664_elements(113) <= OrReduce(convTransposeD_CP_7664_elements(105) & convTransposeD_CP_7664_elements(112));
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_2733/merge_stmt_3167_PhiAck/phi_stmt_3168_ack
      -- 
    phi_stmt_3168_ack_8975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3168_ack_0, ack => convTransposeD_CP_7664_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_2733/merge_stmt_3167_PhiAck/phi_stmt_3174_ack
      -- 
    phi_stmt_3174_ack_8976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3174_ack_0, ack => convTransposeD_CP_7664_elements(115)); -- 
    -- CP-element group 116:  join  fork  transition  place  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: 	70 
    -- CP-element group 116:  members (10) 
      -- CP-element group 116: 	 branch_block_stmt_2733/merge_stmt_3167__exit__
      -- CP-element group 116: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190__entry__
      -- CP-element group 116: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/$entry
      -- CP-element group 116: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_update_start_
      -- CP-element group 116: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_2733/assign_stmt_3185_to_assign_stmt_3190/type_cast_3184_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_2733/merge_stmt_3167_PhiAck/$exit
      -- 
    rr_8652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(116), ack => type_cast_3184_inst_req_0); -- 
    cr_8657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(116), ack => type_cast_3184_inst_req_1); -- 
    convTransposeD_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(114) & convTransposeD_CP_7664_elements(115);
      gj_convTransposeD_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(116), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2965_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2986_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3046_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3077_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2821_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2821_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom65_3088_resized : std_logic_vector(13 downto 0);
    signal R_idxprom65_3088_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_3057_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_3057_scaled : std_logic_vector(13 downto 0);
    signal add21_3028 : std_logic_vector(31 downto 0);
    signal add29_2926 : std_logic_vector(31 downto 0);
    signal add40_2941 : std_logic_vector(31 downto 0);
    signal add55_2998 : std_logic_vector(31 downto 0);
    signal add57_3033 : std_logic_vector(31 downto 0);
    signal add70_3106 : std_logic_vector(31 downto 0);
    signal add_2911 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3058_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3058_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3058_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3058_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3058_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3058_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3089_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3089_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3089_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3089_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3089_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3089_root_address : std_logic_vector(13 downto 0);
    signal arrayidx66_3091 : std_logic_vector(31 downto 0);
    signal arrayidx_3060 : std_logic_vector(31 downto 0);
    signal call_2736 : std_logic_vector(15 downto 0);
    signal cmp81_3142 : std_logic_vector(0 downto 0);
    signal cmp92_3190 : std_logic_vector(0 downto 0);
    signal cmp_3111 : std_logic_vector(0 downto 0);
    signal conv13105_3023 : std_logic_vector(31 downto 0);
    signal conv16_2896 : std_logic_vector(31 downto 0);
    signal conv19_2901 : std_logic_vector(31 downto 0);
    signal conv26_2807 : std_logic_vector(31 downto 0);
    signal conv31_2826 : std_logic_vector(31 downto 0);
    signal conv37_2840 : std_logic_vector(31 downto 0);
    signal conv4_2781 : std_logic_vector(15 downto 0);
    signal conv50_2967 : std_logic_vector(31 downto 0);
    signal conv53_2988 : std_logic_vector(31 downto 0);
    signal conv69_3100 : std_logic_vector(31 downto 0);
    signal conv79_3137 : std_logic_vector(31 downto 0);
    signal conv88_3165 : std_logic_vector(15 downto 0);
    signal conv90_3185 : std_logic_vector(31 downto 0);
    signal conv_2759 : std_logic_vector(15 downto 0);
    signal div3_2777 : std_logic_vector(31 downto 0);
    signal div87_3161 : std_logic_vector(31 downto 0);
    signal div_2755 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2872 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2745 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2767 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2789 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2799 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2815 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2832 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2848 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2860 : std_logic_vector(31 downto 0);
    signal idxprom65_3084 : std_logic_vector(63 downto 0);
    signal idxprom_3053 : std_logic_vector(63 downto 0);
    signal inc85_3155 : std_logic_vector(15 downto 0);
    signal inc_3132 : std_logic_vector(15 downto 0);
    signal indvar_3006 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_3124 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_3174 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2885 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2879 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_3168 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_3019 : std_logic_vector(15 downto 0);
    signal mul20_2916 : std_logic_vector(31 downto 0);
    signal mul27_2921 : std_logic_vector(31 downto 0);
    signal mul38_2936 : std_logic_vector(31 downto 0);
    signal mul54_2993 : std_logic_vector(31 downto 0);
    signal mul56_3003 : std_logic_vector(31 downto 0);
    signal mul_2906 : std_logic_vector(31 downto 0);
    signal ptr_deref_2748_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2748_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2748_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2748_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2748_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2770_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2770_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2770_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2770_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2770_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2792_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2792_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2792_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2792_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2792_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2802_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2802_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2802_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2802_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2802_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2818_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2818_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2818_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2818_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2818_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2835_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2835_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2835_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2835_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2835_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2851_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2851_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2851_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2851_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2851_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2863_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2863_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2863_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2863_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2863_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2875_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2875_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2875_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2875_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2875_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3063_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3063_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3063_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3063_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3063_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3093_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3093_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3093_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3093_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3093_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3093_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext106_2979 : std_logic_vector(31 downto 0);
    signal sext108_3039 : std_logic_vector(31 downto 0);
    signal sext109_3070 : std_logic_vector(31 downto 0);
    signal sext_2958 : std_logic_vector(31 downto 0);
    signal shr64_3079 : std_logic_vector(31 downto 0);
    signal shr_3048 : std_logic_vector(31 downto 0);
    signal sub32_2973 : std_logic_vector(31 downto 0);
    signal sub43_2946 : std_logic_vector(31 downto 0);
    signal sub44_2952 : std_logic_vector(31 downto 0);
    signal sub_2931 : std_logic_vector(31 downto 0);
    signal tmp14_2793 : std_logic_vector(31 downto 0);
    signal tmp25_2803 : std_logic_vector(15 downto 0);
    signal tmp28_2819 : std_logic_vector(31 downto 0);
    signal tmp2_2771 : std_logic_vector(31 downto 0);
    signal tmp30_2822 : std_logic_vector(15 downto 0);
    signal tmp36_2836 : std_logic_vector(15 downto 0);
    signal tmp39_2852 : std_logic_vector(31 downto 0);
    signal tmp48_2864 : std_logic_vector(31 downto 0);
    signal tmp51_2876 : std_logic_vector(31 downto 0);
    signal tmp61_3064 : std_logic_vector(63 downto 0);
    signal tmp_2749 : std_logic_vector(31 downto 0);
    signal type_cast_2753_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2775_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2882_wire : std_logic_vector(15 downto 0);
    signal type_cast_2884_wire : std_logic_vector(15 downto 0);
    signal type_cast_2888_wire : std_logic_vector(15 downto 0);
    signal type_cast_2890_wire : std_logic_vector(15 downto 0);
    signal type_cast_2894_wire : std_logic_vector(31 downto 0);
    signal type_cast_2899_wire : std_logic_vector(31 downto 0);
    signal type_cast_2950_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2956_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2961_wire : std_logic_vector(31 downto 0);
    signal type_cast_2964_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2971_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2977_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2982_wire : std_logic_vector(31 downto 0);
    signal type_cast_2985_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3010_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3012_wire : std_logic_vector(15 downto 0);
    signal type_cast_3017_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3037_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3042_wire : std_logic_vector(31 downto 0);
    signal type_cast_3045_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3051_wire : std_logic_vector(63 downto 0);
    signal type_cast_3068_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3073_wire : std_logic_vector(31 downto 0);
    signal type_cast_3076_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3082_wire : std_logic_vector(63 downto 0);
    signal type_cast_3098_wire : std_logic_vector(31 downto 0);
    signal type_cast_3104_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3122_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3130_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3135_wire : std_logic_vector(31 downto 0);
    signal type_cast_3153_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3159_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3171_wire : std_logic_vector(15 downto 0);
    signal type_cast_3173_wire : std_logic_vector(15 downto 0);
    signal type_cast_3177_wire : std_logic_vector(15 downto 0);
    signal type_cast_3179_wire : std_logic_vector(15 downto 0);
    signal type_cast_3183_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2821_word_address_0 <= "0";
    array_obj_ref_3058_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3058_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3058_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3058_resized_base_address <= "00000000000000";
    array_obj_ref_3089_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3089_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3089_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3089_resized_base_address <= "00000000000000";
    iNsTr_10_2872 <= "00000000000000000000000000000011";
    iNsTr_2_2745 <= "00000000000000000000000000000010";
    iNsTr_3_2767 <= "00000000000000000000000000000011";
    iNsTr_4_2789 <= "00000000000000000000000000000100";
    iNsTr_5_2799 <= "00000000000000000000000000000000";
    iNsTr_6_2815 <= "00000000000000000000000000000011";
    iNsTr_7_2832 <= "00000000000000000000000000000001";
    iNsTr_8_2848 <= "00000000000000000000000000000100";
    iNsTr_9_2860 <= "00000000000000000000000000000100";
    ptr_deref_2748_word_offset_0 <= "0000000";
    ptr_deref_2770_word_offset_0 <= "0000000";
    ptr_deref_2792_word_offset_0 <= "0000000";
    ptr_deref_2802_word_offset_0 <= "0";
    ptr_deref_2818_word_offset_0 <= "0000000";
    ptr_deref_2835_word_offset_0 <= "0";
    ptr_deref_2851_word_offset_0 <= "0000000";
    ptr_deref_2863_word_offset_0 <= "0000000";
    ptr_deref_2875_word_offset_0 <= "0000000";
    ptr_deref_3063_word_offset_0 <= "00000000000000";
    ptr_deref_3093_word_offset_0 <= "00000000000000";
    type_cast_2753_wire_constant <= "00000000000000000000000000000001";
    type_cast_2775_wire_constant <= "00000000000000000000000000000001";
    type_cast_2950_wire_constant <= "00000000000000000000000000010000";
    type_cast_2956_wire_constant <= "11111111111111110000000000000000";
    type_cast_2964_wire_constant <= "00000000000000000000000000010000";
    type_cast_2971_wire_constant <= "00000000000000000000000000010000";
    type_cast_2977_wire_constant <= "11111111111111110000000000000000";
    type_cast_2985_wire_constant <= "00000000000000000000000000010000";
    type_cast_3010_wire_constant <= "0000000000000000";
    type_cast_3017_wire_constant <= "0000000000000100";
    type_cast_3037_wire_constant <= "00000000000000000000000000010000";
    type_cast_3045_wire_constant <= "00000000000000000000000000010010";
    type_cast_3068_wire_constant <= "00000000000000000000000000010000";
    type_cast_3076_wire_constant <= "00000000000000000000000000010010";
    type_cast_3104_wire_constant <= "00000000000000000000000000000100";
    type_cast_3122_wire_constant <= "0000000000000001";
    type_cast_3130_wire_constant <= "0000000000000001";
    type_cast_3153_wire_constant <= "0000000000000001";
    type_cast_3159_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_2879: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2882_wire & type_cast_2884_wire;
      req <= phi_stmt_2879_req_0 & phi_stmt_2879_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2879",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2879_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2879,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2879
    phi_stmt_2885: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2888_wire & type_cast_2890_wire;
      req <= phi_stmt_2885_req_0 & phi_stmt_2885_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2885",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2885_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2885,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2885
    phi_stmt_3006: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3010_wire_constant & type_cast_3012_wire;
      req <= phi_stmt_3006_req_0 & phi_stmt_3006_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3006",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3006_ack_0,
          idata => idata,
          odata => indvar_3006,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3006
    phi_stmt_3168: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3171_wire & type_cast_3173_wire;
      req <= phi_stmt_3168_req_0 & phi_stmt_3168_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3168",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3168_ack_0,
          idata => idata,
          odata => input_dim1x_x2_3168,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3168
    phi_stmt_3174: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3177_wire & type_cast_3179_wire;
      req <= phi_stmt_3174_req_0 & phi_stmt_3174_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3174",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3174_ack_0,
          idata => idata,
          odata => input_dim0x_x0_3174,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3174
    addr_of_3059_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3059_final_reg_req_0;
      addr_of_3059_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3059_final_reg_req_1;
      addr_of_3059_final_reg_ack_1<= rack(0);
      addr_of_3059_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3059_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3058_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_3060,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3090_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3090_final_reg_req_0;
      addr_of_3090_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3090_final_reg_req_1;
      addr_of_3090_final_reg_ack_1<= rack(0);
      addr_of_3090_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3090_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3089_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx66_3091,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2758_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2758_inst_req_0;
      type_cast_2758_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2758_inst_req_1;
      type_cast_2758_inst_ack_1<= rack(0);
      type_cast_2758_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2758_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2755,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2759,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2780_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2780_inst_req_0;
      type_cast_2780_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2780_inst_req_1;
      type_cast_2780_inst_ack_1<= rack(0);
      type_cast_2780_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2780_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div3_2777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_2781,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2806_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2806_inst_req_0;
      type_cast_2806_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2806_inst_req_1;
      type_cast_2806_inst_ack_1<= rack(0);
      type_cast_2806_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2806_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp25_2803,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_2807,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2825_inst_req_0;
      type_cast_2825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2825_inst_req_1;
      type_cast_2825_inst_ack_1<= rack(0);
      type_cast_2825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp30_2822,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_2826,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2839_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2839_inst_req_0;
      type_cast_2839_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2839_inst_req_1;
      type_cast_2839_inst_ack_1<= rack(0);
      type_cast_2839_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2839_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp36_2836,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_2840,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2882_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2882_inst_req_0;
      type_cast_2882_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2882_inst_req_1;
      type_cast_2882_inst_ack_1<= rack(0);
      type_cast_2882_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2882_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_2781,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2882_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2884_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2884_inst_req_0;
      type_cast_2884_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2884_inst_req_1;
      type_cast_2884_inst_ack_1<= rack(0);
      type_cast_2884_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2884_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_3168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2884_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2888_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2888_inst_req_0;
      type_cast_2888_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2888_inst_req_1;
      type_cast_2888_inst_ack_1<= rack(0);
      type_cast_2888_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2888_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2759,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2888_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2890_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2890_inst_req_0;
      type_cast_2890_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2890_inst_req_1;
      type_cast_2890_inst_ack_1<= rack(0);
      type_cast_2890_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2890_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_3174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2890_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2895_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2895_inst_req_0;
      type_cast_2895_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2895_inst_req_1;
      type_cast_2895_inst_ack_1<= rack(0);
      type_cast_2895_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2895_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2894_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_2896,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2900_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2900_inst_req_0;
      type_cast_2900_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2900_inst_req_1;
      type_cast_2900_inst_ack_1<= rack(0);
      type_cast_2900_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2900_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2899_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_2901,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2961_inst
    process(sext_2958) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2958(31 downto 0);
      type_cast_2961_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2966_inst
    process(ASHR_i32_i32_2965_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2965_wire(31 downto 0);
      conv50_2967 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2982_inst
    process(sext106_2979) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext106_2979(31 downto 0);
      type_cast_2982_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2987_inst
    process(ASHR_i32_i32_2986_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2986_wire(31 downto 0);
      conv53_2988 <= tmp_var; -- 
    end process;
    type_cast_3012_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3012_inst_req_0;
      type_cast_3012_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3012_inst_req_1;
      type_cast_3012_inst_ack_1<= rack(0);
      type_cast_3012_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3012_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_3124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3012_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3022_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3022_inst_req_0;
      type_cast_3022_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3022_inst_req_1;
      type_cast_3022_inst_ack_1<= rack(0);
      type_cast_3022_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3022_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_3019,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13105_3023,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3042_inst
    process(sext108_3039) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext108_3039(31 downto 0);
      type_cast_3042_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3047_inst
    process(ASHR_i32_i32_3046_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3046_wire(31 downto 0);
      shr_3048 <= tmp_var; -- 
    end process;
    type_cast_3052_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3052_inst_req_0;
      type_cast_3052_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3052_inst_req_1;
      type_cast_3052_inst_ack_1<= rack(0);
      type_cast_3052_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3052_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3051_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_3053,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3073_inst
    process(sext109_3070) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext109_3070(31 downto 0);
      type_cast_3073_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3078_inst
    process(ASHR_i32_i32_3077_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3077_wire(31 downto 0);
      shr64_3079 <= tmp_var; -- 
    end process;
    type_cast_3083_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3083_inst_req_0;
      type_cast_3083_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3083_inst_req_1;
      type_cast_3083_inst_ack_1<= rack(0);
      type_cast_3083_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3083_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3082_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom65_3084,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3099_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3099_inst_req_0;
      type_cast_3099_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3099_inst_req_1;
      type_cast_3099_inst_ack_1<= rack(0);
      type_cast_3099_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3099_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3098_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_3100,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3136_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3136_inst_req_0;
      type_cast_3136_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3136_inst_req_1;
      type_cast_3136_inst_ack_1<= rack(0);
      type_cast_3136_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3136_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3135_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_3137,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3164_inst_req_0;
      type_cast_3164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3164_inst_req_1;
      type_cast_3164_inst_ack_1<= rack(0);
      type_cast_3164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div87_3161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_3165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3171_inst_req_0;
      type_cast_3171_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3171_inst_req_1;
      type_cast_3171_inst_ack_1<= rack(0);
      type_cast_3171_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3171_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv88_3165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3171_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3173_inst_req_0;
      type_cast_3173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3173_inst_req_1;
      type_cast_3173_inst_ack_1<= rack(0);
      type_cast_3173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_3132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3173_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3177_inst_req_0;
      type_cast_3177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3177_inst_req_1;
      type_cast_3177_inst_ack_1<= rack(0);
      type_cast_3177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc85_3155,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3177_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3179_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3179_inst_req_0;
      type_cast_3179_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3179_inst_req_1;
      type_cast_3179_inst_ack_1<= rack(0);
      type_cast_3179_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3179_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2x_xph_2885,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3179_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3184_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3184_inst_req_0;
      type_cast_3184_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3184_inst_req_1;
      type_cast_3184_inst_ack_1<= rack(0);
      type_cast_3184_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3184_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3183_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_3185,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2821_gather_scatter
    process(LOAD_padding_2821_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2821_data_0;
      ov(15 downto 0) := iv;
      tmp30_2822 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3058_index_1_rename
    process(R_idxprom_3057_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_3057_resized;
      ov(13 downto 0) := iv;
      R_idxprom_3057_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3058_index_1_resize
    process(idxprom_3053) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_3053;
      ov := iv(13 downto 0);
      R_idxprom_3057_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3058_root_address_inst
    process(array_obj_ref_3058_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3058_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3058_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3089_index_1_rename
    process(R_idxprom65_3088_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom65_3088_resized;
      ov(13 downto 0) := iv;
      R_idxprom65_3088_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3089_index_1_resize
    process(idxprom65_3084) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom65_3084;
      ov := iv(13 downto 0);
      R_idxprom65_3088_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3089_root_address_inst
    process(array_obj_ref_3089_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3089_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3089_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2748_addr_0
    process(ptr_deref_2748_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2748_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2748_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2748_base_resize
    process(iNsTr_2_2745) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2745;
      ov := iv(6 downto 0);
      ptr_deref_2748_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2748_gather_scatter
    process(ptr_deref_2748_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2748_data_0;
      ov(31 downto 0) := iv;
      tmp_2749 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2748_root_address_inst
    process(ptr_deref_2748_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2748_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2748_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2770_addr_0
    process(ptr_deref_2770_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2770_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2770_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2770_base_resize
    process(iNsTr_3_2767) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2767;
      ov := iv(6 downto 0);
      ptr_deref_2770_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2770_gather_scatter
    process(ptr_deref_2770_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2770_data_0;
      ov(31 downto 0) := iv;
      tmp2_2771 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2770_root_address_inst
    process(ptr_deref_2770_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2770_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2770_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2792_addr_0
    process(ptr_deref_2792_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2792_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2792_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2792_base_resize
    process(iNsTr_4_2789) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2789;
      ov := iv(6 downto 0);
      ptr_deref_2792_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2792_gather_scatter
    process(ptr_deref_2792_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2792_data_0;
      ov(31 downto 0) := iv;
      tmp14_2793 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2792_root_address_inst
    process(ptr_deref_2792_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2792_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2792_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2802_addr_0
    process(ptr_deref_2802_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2802_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2802_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2802_base_resize
    process(iNsTr_5_2799) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2799;
      ov := iv(0 downto 0);
      ptr_deref_2802_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2802_gather_scatter
    process(ptr_deref_2802_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2802_data_0;
      ov(15 downto 0) := iv;
      tmp25_2803 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2802_root_address_inst
    process(ptr_deref_2802_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2802_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2802_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2818_addr_0
    process(ptr_deref_2818_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2818_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2818_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2818_base_resize
    process(iNsTr_6_2815) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2815;
      ov := iv(6 downto 0);
      ptr_deref_2818_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2818_gather_scatter
    process(ptr_deref_2818_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2818_data_0;
      ov(31 downto 0) := iv;
      tmp28_2819 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2818_root_address_inst
    process(ptr_deref_2818_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2818_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2818_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2835_addr_0
    process(ptr_deref_2835_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2835_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2835_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2835_base_resize
    process(iNsTr_7_2832) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2832;
      ov := iv(0 downto 0);
      ptr_deref_2835_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2835_gather_scatter
    process(ptr_deref_2835_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2835_data_0;
      ov(15 downto 0) := iv;
      tmp36_2836 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2835_root_address_inst
    process(ptr_deref_2835_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2835_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2835_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2851_addr_0
    process(ptr_deref_2851_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2851_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2851_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2851_base_resize
    process(iNsTr_8_2848) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2848;
      ov := iv(6 downto 0);
      ptr_deref_2851_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2851_gather_scatter
    process(ptr_deref_2851_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2851_data_0;
      ov(31 downto 0) := iv;
      tmp39_2852 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2851_root_address_inst
    process(ptr_deref_2851_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2851_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2851_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2863_addr_0
    process(ptr_deref_2863_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2863_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2863_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2863_base_resize
    process(iNsTr_9_2860) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2860;
      ov := iv(6 downto 0);
      ptr_deref_2863_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2863_gather_scatter
    process(ptr_deref_2863_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2863_data_0;
      ov(31 downto 0) := iv;
      tmp48_2864 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2863_root_address_inst
    process(ptr_deref_2863_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2863_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2863_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2875_addr_0
    process(ptr_deref_2875_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2875_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2875_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2875_base_resize
    process(iNsTr_10_2872) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2872;
      ov := iv(6 downto 0);
      ptr_deref_2875_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2875_gather_scatter
    process(ptr_deref_2875_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2875_data_0;
      ov(31 downto 0) := iv;
      tmp51_2876 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2875_root_address_inst
    process(ptr_deref_2875_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2875_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2875_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3063_addr_0
    process(ptr_deref_3063_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3063_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3063_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3063_base_resize
    process(arrayidx_3060) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_3060;
      ov := iv(13 downto 0);
      ptr_deref_3063_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3063_gather_scatter
    process(ptr_deref_3063_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3063_data_0;
      ov(63 downto 0) := iv;
      tmp61_3064 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3063_root_address_inst
    process(ptr_deref_3063_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3063_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3063_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3093_addr_0
    process(ptr_deref_3093_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3093_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3093_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3093_base_resize
    process(arrayidx66_3091) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx66_3091;
      ov := iv(13 downto 0);
      ptr_deref_3093_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3093_gather_scatter
    process(tmp61_3064) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp61_3064;
      ov(63 downto 0) := iv;
      ptr_deref_3093_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3093_root_address_inst
    process(ptr_deref_3093_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3093_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3093_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_3112_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_3111;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3112_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3112_branch_req_0,
          ack0 => if_stmt_3112_branch_ack_0,
          ack1 => if_stmt_3112_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3143_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp81_3142;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3143_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3143_branch_req_0,
          ack0 => if_stmt_3143_branch_ack_0,
          ack1 => if_stmt_3143_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3191_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp92_3190;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3191_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3191_branch_req_0,
          ack0 => if_stmt_3191_branch_ack_0,
          ack1 => if_stmt_3191_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3123_inst
    process(indvar_3006) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_3006, type_cast_3122_wire_constant, tmp_var);
      indvarx_xnext_3124 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3131_inst
    process(input_dim1x_x1x_xph_2879) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2879, type_cast_3130_wire_constant, tmp_var);
      inc_3132 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3154_inst
    process(input_dim0x_x2x_xph_2885) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_2885, type_cast_3153_wire_constant, tmp_var);
      inc85_3155 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2910_inst
    process(mul_2906, conv16_2896) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2906, conv16_2896, tmp_var);
      add_2911 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2925_inst
    process(mul27_2921, tmp28_2819) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul27_2921, tmp28_2819, tmp_var);
      add29_2926 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2940_inst
    process(mul38_2936, tmp39_2852) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul38_2936, tmp39_2852, tmp_var);
      add40_2941 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2957_inst
    process(sub44_2952) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub44_2952, type_cast_2956_wire_constant, tmp_var);
      sext_2958 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2978_inst
    process(sub32_2973) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub32_2973, type_cast_2977_wire_constant, tmp_var);
      sext106_2979 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2997_inst
    process(conv50_2967, mul54_2993) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv50_2967, mul54_2993, tmp_var);
      add55_2998 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3027_inst
    process(mul20_2916, conv13105_3023) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul20_2916, conv13105_3023, tmp_var);
      add21_3028 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3032_inst
    process(mul56_3003, conv13105_3023) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul56_3003, conv13105_3023, tmp_var);
      add57_3033 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3105_inst
    process(conv69_3100) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv69_3100, type_cast_3104_wire_constant, tmp_var);
      add70_3106 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2965_inst
    process(type_cast_2961_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2961_wire, type_cast_2964_wire_constant, tmp_var);
      ASHR_i32_i32_2965_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2986_inst
    process(type_cast_2982_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2982_wire, type_cast_2985_wire_constant, tmp_var);
      ASHR_i32_i32_2986_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3046_inst
    process(type_cast_3042_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3042_wire, type_cast_3045_wire_constant, tmp_var);
      ASHR_i32_i32_3046_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3077_inst
    process(type_cast_3073_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3073_wire, type_cast_3076_wire_constant, tmp_var);
      ASHR_i32_i32_3077_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3141_inst
    process(conv79_3137, tmp2_2771) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv79_3137, tmp2_2771, tmp_var);
      cmp81_3142 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3189_inst
    process(conv90_3185, tmp_2749) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv90_3185, tmp_2749, tmp_var);
      cmp92_3190 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2754_inst
    process(tmp_2749) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2749, type_cast_2753_wire_constant, tmp_var);
      div_2755 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2776_inst
    process(tmp2_2771) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2771, type_cast_2775_wire_constant, tmp_var);
      div3_2777 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3160_inst
    process(tmp2_2771) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2771, type_cast_3159_wire_constant, tmp_var);
      div87_3161 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3018_inst
    process(indvar_3006) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_3006, type_cast_3017_wire_constant, tmp_var);
      input_dim2x_x1_3019 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2905_inst
    process(tmp2_2771, conv19_2901) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_2771, conv19_2901, tmp_var);
      mul_2906 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2915_inst
    process(add_2911, tmp14_2793) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2911, tmp14_2793, tmp_var);
      mul20_2916 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2920_inst
    process(conv26_2807, conv19_2901) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv26_2807, conv19_2901, tmp_var);
      mul27_2921 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2935_inst
    process(conv37_2840, conv16_2896) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv37_2840, conv16_2896, tmp_var);
      mul38_2936 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2992_inst
    process(tmp51_2876, conv53_2988) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp51_2876, conv53_2988, tmp_var);
      mul54_2993 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3002_inst
    process(add55_2998, tmp48_2864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add55_2998, tmp48_2864, tmp_var);
      mul56_3003 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2951_inst
    process(sub43_2946) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub43_2946, type_cast_2950_wire_constant, tmp_var);
      sub44_2952 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2972_inst
    process(sub_2931) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2931, type_cast_2971_wire_constant, tmp_var);
      sub32_2973 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3038_inst
    process(add21_3028) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add21_3028, type_cast_3037_wire_constant, tmp_var);
      sext108_3039 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3069_inst
    process(add57_3033) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add57_3033, type_cast_3068_wire_constant, tmp_var);
      sext109_3070 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2930_inst
    process(add29_2926, conv31_2826) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add29_2926, conv31_2826, tmp_var);
      sub_2931 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2945_inst
    process(add40_2941, conv31_2826) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add40_2941, conv31_2826, tmp_var);
      sub43_2946 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_3110_inst
    process(add70_3106, tmp14_2793) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add70_3106, tmp14_2793, tmp_var);
      cmp_3111 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_3058_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_3057_scaled;
      array_obj_ref_3058_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3058_index_offset_req_0;
      array_obj_ref_3058_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3058_index_offset_req_1;
      array_obj_ref_3058_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_3089_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom65_3088_scaled;
      array_obj_ref_3089_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3089_index_offset_req_0;
      array_obj_ref_3089_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3089_index_offset_req_1;
      array_obj_ref_3089_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- unary operator type_cast_2894_inst
    process(input_dim1x_x1x_xph_2879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_2879, tmp_var);
      type_cast_2894_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2899_inst
    process(input_dim0x_x2x_xph_2885) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_2885, tmp_var);
      type_cast_2899_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3051_inst
    process(shr_3048) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_3048, tmp_var);
      type_cast_3051_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3082_inst
    process(shr64_3079) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr64_3079, tmp_var);
      type_cast_3082_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3098_inst
    process(input_dim2x_x1_3019) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_3019, tmp_var);
      type_cast_3098_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3135_inst
    process(inc_3132) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_3132, tmp_var);
      type_cast_3135_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3183_inst
    process(input_dim0x_x0_3174) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_3174, tmp_var);
      type_cast_3183_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2821_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2821_load_0_req_0;
      LOAD_padding_2821_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2821_load_0_req_1;
      LOAD_padding_2821_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2821_word_address_0;
      LOAD_padding_2821_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2748_load_0 ptr_deref_2770_load_0 ptr_deref_2792_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2748_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2770_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2792_load_0_req_0;
      ptr_deref_2748_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2770_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2792_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2748_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2770_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2792_load_0_req_1;
      ptr_deref_2748_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2770_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2792_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2748_word_address_0 & ptr_deref_2770_word_address_0 & ptr_deref_2792_word_address_0;
      ptr_deref_2748_data_0 <= data_out(95 downto 64);
      ptr_deref_2770_data_0 <= data_out(63 downto 32);
      ptr_deref_2792_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2835_load_0 ptr_deref_2802_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2835_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2802_load_0_req_0;
      ptr_deref_2835_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2802_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2835_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2802_load_0_req_1;
      ptr_deref_2835_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2802_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2835_word_address_0 & ptr_deref_2802_word_address_0;
      ptr_deref_2835_data_0 <= data_out(31 downto 16);
      ptr_deref_2802_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(15 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2818_load_0 ptr_deref_2851_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2818_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2851_load_0_req_0;
      ptr_deref_2818_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2851_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2818_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2851_load_0_req_1;
      ptr_deref_2818_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2851_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2818_word_address_0 & ptr_deref_2851_word_address_0;
      ptr_deref_2818_data_0 <= data_out(63 downto 32);
      ptr_deref_2851_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2875_load_0 ptr_deref_2863_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2875_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2863_load_0_req_0;
      ptr_deref_2875_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2863_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2875_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2863_load_0_req_1;
      ptr_deref_2875_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2863_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2875_word_address_0 & ptr_deref_2863_word_address_0;
      ptr_deref_2875_data_0 <= data_out(63 downto 32);
      ptr_deref_2863_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_3063_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3063_load_0_req_0;
      ptr_deref_3063_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3063_load_0_req_1;
      ptr_deref_3063_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3063_word_address_0;
      ptr_deref_3063_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_3093_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3093_store_0_req_0;
      ptr_deref_3093_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3093_store_0_req_1;
      ptr_deref_3093_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3093_word_address_0;
      data_in <= ptr_deref_3093_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2735_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_start_2735_inst_req_0;
      RPIPE_Block3_start_2735_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_start_2735_inst_req_1;
      RPIPE_Block3_start_2735_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2736 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_3199_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_3199_inst_req_0;
      WPIPE_Block3_done_3199_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_3199_inst_req_1;
      WPIPE_Block3_done_3199_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2736;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_3266_start: Boolean;
  signal sendOutput_CP_3266_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal addr_of_1201_final_reg_req_0 : boolean;
  signal addr_of_1201_final_reg_ack_0 : boolean;
  signal if_stmt_1144_branch_ack_0 : boolean;
  signal ptr_deref_1102_load_0_req_1 : boolean;
  signal ptr_deref_1102_load_0_ack_1 : boolean;
  signal ptr_deref_1102_load_0_ack_0 : boolean;
  signal ptr_deref_1205_load_0_req_0 : boolean;
  signal ptr_deref_1102_load_0_req_0 : boolean;
  signal array_obj_ref_1200_index_offset_ack_1 : boolean;
  signal array_obj_ref_1200_index_offset_req_1 : boolean;
  signal ptr_deref_1114_load_0_ack_1 : boolean;
  signal ptr_deref_1205_load_0_req_1 : boolean;
  signal ptr_deref_1114_load_0_req_1 : boolean;
  signal array_obj_ref_1200_index_offset_ack_0 : boolean;
  signal type_cast_1229_inst_req_1 : boolean;
  signal type_cast_1219_inst_req_0 : boolean;
  signal type_cast_1209_inst_req_1 : boolean;
  signal type_cast_1239_inst_req_1 : boolean;
  signal type_cast_1209_inst_ack_1 : boolean;
  signal type_cast_1229_inst_req_0 : boolean;
  signal ptr_deref_1205_load_0_ack_1 : boolean;
  signal type_cast_1229_inst_ack_0 : boolean;
  signal type_cast_1219_inst_ack_0 : boolean;
  signal type_cast_1239_inst_ack_1 : boolean;
  signal ptr_deref_1205_load_0_ack_0 : boolean;
  signal addr_of_1201_final_reg_req_1 : boolean;
  signal type_cast_1229_inst_ack_1 : boolean;
  signal addr_of_1201_final_reg_ack_1 : boolean;
  signal ptr_deref_1126_load_0_ack_0 : boolean;
  signal ptr_deref_1126_load_0_req_0 : boolean;
  signal type_cast_1269_inst_ack_1 : boolean;
  signal type_cast_1249_inst_req_0 : boolean;
  signal type_cast_1249_inst_ack_0 : boolean;
  signal if_stmt_1144_branch_req_0 : boolean;
  signal type_cast_1279_inst_req_1 : boolean;
  signal type_cast_1279_inst_ack_1 : boolean;
  signal type_cast_1239_inst_req_0 : boolean;
  signal type_cast_1209_inst_req_0 : boolean;
  signal type_cast_1269_inst_req_0 : boolean;
  signal type_cast_1269_inst_ack_0 : boolean;
  signal ptr_deref_1114_load_0_req_0 : boolean;
  signal type_cast_1249_inst_req_1 : boolean;
  signal type_cast_1249_inst_ack_1 : boolean;
  signal ptr_deref_1126_load_0_req_1 : boolean;
  signal type_cast_1219_inst_req_1 : boolean;
  signal ptr_deref_1114_load_0_ack_0 : boolean;
  signal type_cast_1209_inst_ack_0 : boolean;
  signal ptr_deref_1126_load_0_ack_1 : boolean;
  signal type_cast_1269_inst_req_1 : boolean;
  signal type_cast_1239_inst_ack_0 : boolean;
  signal type_cast_1279_inst_req_0 : boolean;
  signal type_cast_1279_inst_ack_0 : boolean;
  signal type_cast_1219_inst_ack_1 : boolean;
  signal type_cast_1171_inst_ack_0 : boolean;
  signal type_cast_1171_inst_req_0 : boolean;
  signal type_cast_1259_inst_req_0 : boolean;
  signal type_cast_1259_inst_ack_0 : boolean;
  signal type_cast_1171_inst_ack_1 : boolean;
  signal array_obj_ref_1200_index_offset_req_0 : boolean;
  signal type_cast_1259_inst_req_1 : boolean;
  signal type_cast_1171_inst_req_1 : boolean;
  signal type_cast_1259_inst_ack_1 : boolean;
  signal if_stmt_1144_branch_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1 : boolean;
  signal if_stmt_1316_branch_req_0 : boolean;
  signal if_stmt_1316_branch_ack_1 : boolean;
  signal if_stmt_1316_branch_ack_0 : boolean;
  signal phi_stmt_1188_req_0 : boolean;
  signal type_cast_1194_inst_req_0 : boolean;
  signal type_cast_1194_inst_ack_0 : boolean;
  signal type_cast_1194_inst_req_1 : boolean;
  signal type_cast_1194_inst_ack_1 : boolean;
  signal phi_stmt_1188_req_1 : boolean;
  signal phi_stmt_1188_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_3266_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_3266_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_3266_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_3266_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_3266: Block -- control-path 
    signal sendOutput_CP_3266_elements: BooleanArray(66 downto 0);
    -- 
  begin -- 
    sendOutput_CP_3266_elements(0) <= sendOutput_CP_3266_start;
    sendOutput_CP_3266_symbol <= sendOutput_CP_3266_elements(66);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (83) 
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143__entry__
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1091/branch_block_stmt_1091__entry__
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1091/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_root_address_calculated
      -- 
    cr_3340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1102_load_0_req_1); -- 
    rr_3329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1102_load_0_req_0); -- 
    cr_3390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1114_load_0_req_1); -- 
    rr_3429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1126_load_0_req_0); -- 
    rr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1114_load_0_req_0); -- 
    cr_3440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1126_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Sample/word_access_start/$exit
      -- 
    ra_3330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1102_load_0_ack_0, ack => sendOutput_CP_3266_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/ptr_deref_1102_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/ptr_deref_1102_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/ptr_deref_1102_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1102_Update/ptr_deref_1102_Merge/merge_ack
      -- 
    ca_3341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1102_load_0_ack_1, ack => sendOutput_CP_3266_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Sample/word_access_start/word_0/ra
      -- 
    ra_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1114_load_0_ack_0, ack => sendOutput_CP_3266_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/ptr_deref_1114_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/ptr_deref_1114_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/ptr_deref_1114_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/ptr_deref_1114_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1114_Update/word_access_complete/$exit
      -- 
    ca_3391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1114_load_0_ack_1, ack => sendOutput_CP_3266_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_sample_completed_
      -- 
    ra_3430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1126_load_0_ack_0, ack => sendOutput_CP_3266_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/ptr_deref_1126_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/ptr_deref_1126_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/ptr_deref_1126_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/ptr_deref_1126_Update/ptr_deref_1126_Merge/$entry
      -- 
    ca_3441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1126_load_0_ack_1, ack => sendOutput_CP_3266_elements(6)); -- 
    -- CP-element group 7:  branch  join  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (10) 
      -- CP-element group 7: 	 branch_block_stmt_1091/if_stmt_1144_eval_test/$entry
      -- CP-element group 7: 	 branch_block_stmt_1091/if_stmt_1144__entry__
      -- CP-element group 7: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143__exit__
      -- CP-element group 7: 	 branch_block_stmt_1091/if_stmt_1144_dead_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_1091/assign_stmt_1099_to_assign_stmt_1143/$exit
      -- CP-element group 7: 	 branch_block_stmt_1091/if_stmt_1144_eval_test/$exit
      -- CP-element group 7: 	 branch_block_stmt_1091/if_stmt_1144_eval_test/branch_req
      -- CP-element group 7: 	 branch_block_stmt_1091/R_cmp73_1145_place
      -- CP-element group 7: 	 branch_block_stmt_1091/if_stmt_1144_if_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_1091/if_stmt_1144_else_link/$entry
      -- 
    branch_req_3454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(7), ack => if_stmt_1144_branch_req_0); -- 
    sendOutput_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "sendOutput_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(6) & sendOutput_CP_3266_elements(4) & sendOutput_CP_3266_elements(2);
      gj_sendOutput_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (18) 
      -- CP-element group 8: 	 branch_block_stmt_1091/if_stmt_1144_if_link/$exit
      -- CP-element group 8: 	 branch_block_stmt_1091/entry_bbx_xnph
      -- CP-element group 8: 	 branch_block_stmt_1091/merge_stmt_1150__exit__
      -- CP-element group 8: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185__entry__
      -- CP-element group 8: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/$entry
      -- CP-element group 8: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1091/if_stmt_1144_if_link/if_choice_transition
      -- CP-element group 8: 	 branch_block_stmt_1091/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_1091/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 8: 	 branch_block_stmt_1091/merge_stmt_1150_PhiReqMerge
      -- CP-element group 8: 	 branch_block_stmt_1091/merge_stmt_1150_PhiAck/$entry
      -- CP-element group 8: 	 branch_block_stmt_1091/merge_stmt_1150_PhiAck/$exit
      -- CP-element group 8: 	 branch_block_stmt_1091/merge_stmt_1150_PhiAck/dummy
      -- 
    if_choice_transition_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1144_branch_ack_1, ack => sendOutput_CP_3266_elements(8)); -- 
    rr_3476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(8), ack => type_cast_1171_inst_req_0); -- 
    cr_3481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(8), ack => type_cast_1171_inst_req_1); -- 
    -- CP-element group 9:  transition  place  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	66 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1091/if_stmt_1144_else_link/else_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_1091/entry_forx_xend
      -- CP-element group 9: 	 branch_block_stmt_1091/if_stmt_1144_else_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_1091/entry_forx_xend_PhiReq/$entry
      -- CP-element group 9: 	 branch_block_stmt_1091/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_3463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1144_branch_ack_0, ack => sendOutput_CP_3266_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_sample_completed_
      -- 
    ra_3477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_0, ack => sendOutput_CP_3266_elements(10)); -- 
    -- CP-element group 11:  transition  place  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	60 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185__exit__
      -- CP-element group 11: 	 branch_block_stmt_1091/bbx_xnph_forx_xbody
      -- CP-element group 11: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/$exit
      -- CP-element group 11: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1091/assign_stmt_1156_to_assign_stmt_1185/type_cast_1171_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1091/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 11: 	 branch_block_stmt_1091/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1188/$entry
      -- CP-element group 11: 	 branch_block_stmt_1091/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/$entry
      -- 
    ca_3482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_1, ack => sendOutput_CP_3266_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	65 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	57 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_final_index_sum_regn_sample_complete
      -- CP-element group 12: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_final_index_sum_regn_Sample/ack
      -- CP-element group 12: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_final_index_sum_regn_Sample/$exit
      -- 
    ack_3511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1200_index_offset_ack_0, ack => sendOutput_CP_3266_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	65 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (11) 
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_request/$entry
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_offset_calculated
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_request/req
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_final_index_sum_regn_Update/ack
      -- CP-element group 13: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_final_index_sum_regn_Update/$exit
      -- 
    ack_3516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1200_index_offset_ack_1, ack => sendOutput_CP_3266_elements(13)); -- 
    req_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(13), ack => addr_of_1201_final_reg_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_request/$exit
      -- CP-element group 14: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_request/ack
      -- CP-element group 14: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_sample_completed_
      -- 
    ack_3526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1201_final_reg_ack_0, ack => sendOutput_CP_3266_elements(14)); -- 
    -- CP-element group 15:  join  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	65 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (24) 
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_base_addr_resize/$exit
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_base_addr_resize/$entry
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_base_address_resized
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Sample/word_access_start/word_0/rr
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_base_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Sample/word_access_start/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_complete/ack
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_base_addr_resize/base_resize_req
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_base_addr_resize/base_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Sample/word_access_start/$entry
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_base_plus_offset/sum_rename_req
      -- 
    ack_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1201_final_reg_ack_1, ack => sendOutput_CP_3266_elements(15)); -- 
    rr_3564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(15), ack => ptr_deref_1205_load_0_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Sample/word_access_start/word_0/ra
      -- CP-element group 16: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Sample/word_access_start/$exit
      -- 
    ra_3565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1205_load_0_ack_0, ack => sendOutput_CP_3266_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	65 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: 	24 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	32 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	28 
    -- CP-element group 17: 	26 
    -- CP-element group 17:  members (33) 
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/ptr_deref_1205_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/ptr_deref_1205_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/ptr_deref_1205_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/ptr_deref_1205_Merge/merge_ack
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_sample_start_
      -- 
    ca_3576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1205_load_0_ack_1, ack => sendOutput_CP_3266_elements(17)); -- 
    rr_3631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1239_inst_req_0); -- 
    rr_3589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1209_inst_req_0); -- 
    rr_3603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1219_inst_req_0); -- 
    rr_3687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1279_inst_req_0); -- 
    rr_3617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1229_inst_req_0); -- 
    rr_3659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1259_inst_req_0); -- 
    rr_3673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1269_inst_req_0); -- 
    rr_3645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1249_inst_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_Sample/ra
      -- 
    ra_3590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1209_inst_ack_0, ack => sendOutput_CP_3266_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	65 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	54 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_update_completed_
      -- 
    ca_3595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1209_inst_ack_1, ack => sendOutput_CP_3266_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_Sample/$exit
      -- 
    ra_3604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1219_inst_ack_0, ack => sendOutput_CP_3266_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	65 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	51 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_Update/ca
      -- 
    ca_3609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1219_inst_ack_1, ack => sendOutput_CP_3266_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	17 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_Sample/$exit
      -- 
    ra_3618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1229_inst_ack_0, ack => sendOutput_CP_3266_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	65 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	48 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_update_completed_
      -- 
    ca_3623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1229_inst_ack_1, ack => sendOutput_CP_3266_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	17 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_Sample/ra
      -- 
    ra_3632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1239_inst_ack_0, ack => sendOutput_CP_3266_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	65 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	45 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_update_completed_
      -- 
    ca_3637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1239_inst_ack_1, ack => sendOutput_CP_3266_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	17 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_sample_completed_
      -- 
    ra_3646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1249_inst_ack_0, ack => sendOutput_CP_3266_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	65 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	42 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_Update/ca
      -- 
    ca_3651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1249_inst_ack_1, ack => sendOutput_CP_3266_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	17 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_Sample/ra
      -- 
    ra_3660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1259_inst_ack_0, ack => sendOutput_CP_3266_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	65 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	39 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_Update/ca
      -- 
    ca_3665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1259_inst_ack_1, ack => sendOutput_CP_3266_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_sample_completed_
      -- 
    ra_3674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1269_inst_ack_0, ack => sendOutput_CP_3266_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	65 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	36 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_Update/$exit
      -- 
    ca_3679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1269_inst_ack_1, ack => sendOutput_CP_3266_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_Sample/ra
      -- 
    ra_3688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_0, ack => sendOutput_CP_3266_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	65 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_Sample/req
      -- 
    ca_3693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_1, ack => sendOutput_CP_3266_elements(33)); -- 
    req_3701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(33), ack => WPIPE_ConvTranspose_output_pipe_1281_inst_req_0); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_Update/req
      -- 
    ack_3702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0, ack => sendOutput_CP_3266_elements(34)); -- 
    req_3706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(34), ack => WPIPE_ConvTranspose_output_pipe_1281_inst_req_1); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1281_Update/ack
      -- 
    ack_3707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1, ack => sendOutput_CP_3266_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: 	31 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_Sample/req
      -- 
    req_3715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(36), ack => WPIPE_ConvTranspose_output_pipe_1284_inst_req_0); -- 
    sendOutput_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(35) & sendOutput_CP_3266_elements(31);
      gj_sendOutput_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_Sample/ack
      -- CP-element group 37: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_Update/req
      -- 
    ack_3716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0, ack => sendOutput_CP_3266_elements(37)); -- 
    req_3720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(37), ack => WPIPE_ConvTranspose_output_pipe_1284_inst_req_1); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1284_Update/ack
      -- 
    ack_3721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1, ack => sendOutput_CP_3266_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: 	29 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_Sample/req
      -- 
    req_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(39), ack => WPIPE_ConvTranspose_output_pipe_1287_inst_req_0); -- 
    sendOutput_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(38) & sendOutput_CP_3266_elements(29);
      gj_sendOutput_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_update_start_
      -- CP-element group 40: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_Update/req
      -- 
    ack_3730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0, ack => sendOutput_CP_3266_elements(40)); -- 
    req_3734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(40), ack => WPIPE_ConvTranspose_output_pipe_1287_inst_req_1); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1287_Update/ack
      -- 
    ack_3735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1, ack => sendOutput_CP_3266_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	27 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_Sample/req
      -- 
    req_3743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(42), ack => WPIPE_ConvTranspose_output_pipe_1290_inst_req_0); -- 
    sendOutput_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(41) & sendOutput_CP_3266_elements(27);
      gj_sendOutput_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_Update/req
      -- 
    ack_3744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0, ack => sendOutput_CP_3266_elements(43)); -- 
    req_3748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(43), ack => WPIPE_ConvTranspose_output_pipe_1290_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1290_Update/ack
      -- 
    ack_3749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1, ack => sendOutput_CP_3266_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	25 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_Sample/req
      -- 
    req_3757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(45), ack => WPIPE_ConvTranspose_output_pipe_1293_inst_req_0); -- 
    sendOutput_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(44) & sendOutput_CP_3266_elements(25);
      gj_sendOutput_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_Update/req
      -- 
    ack_3758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0, ack => sendOutput_CP_3266_elements(46)); -- 
    req_3762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(46), ack => WPIPE_ConvTranspose_output_pipe_1293_inst_req_1); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1293_Update/ack
      -- 
    ack_3763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1, ack => sendOutput_CP_3266_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	23 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_Sample/req
      -- 
    req_3771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(48), ack => WPIPE_ConvTranspose_output_pipe_1296_inst_req_0); -- 
    sendOutput_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(23) & sendOutput_CP_3266_elements(47);
      gj_sendOutput_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_Update/req
      -- 
    ack_3772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0, ack => sendOutput_CP_3266_elements(49)); -- 
    req_3776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(49), ack => WPIPE_ConvTranspose_output_pipe_1296_inst_req_1); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1296_Update/ack
      -- 
    ack_3777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1, ack => sendOutput_CP_3266_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: 	21 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_Sample/req
      -- 
    req_3785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(51), ack => WPIPE_ConvTranspose_output_pipe_1299_inst_req_0); -- 
    sendOutput_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(50) & sendOutput_CP_3266_elements(21);
      gj_sendOutput_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_Update/req
      -- 
    ack_3786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0, ack => sendOutput_CP_3266_elements(52)); -- 
    req_3790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(52), ack => WPIPE_ConvTranspose_output_pipe_1299_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1299_Update/ack
      -- 
    ack_3791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1, ack => sendOutput_CP_3266_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	19 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_Sample/req
      -- 
    req_3799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(54), ack => WPIPE_ConvTranspose_output_pipe_1302_inst_req_0); -- 
    sendOutput_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(19) & sendOutput_CP_3266_elements(53);
      gj_sendOutput_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_Update/req
      -- 
    ack_3800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0, ack => sendOutput_CP_3266_elements(55)); -- 
    req_3804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(55), ack => WPIPE_ConvTranspose_output_pipe_1302_inst_req_1); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/WPIPE_ConvTranspose_output_pipe_1302_Update/ack
      -- 
    ack_3805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1, ack => sendOutput_CP_3266_elements(56)); -- 
    -- CP-element group 57:  branch  join  transition  place  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	12 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (10) 
      -- CP-element group 57: 	 branch_block_stmt_1091/if_stmt_1316__entry__
      -- CP-element group 57: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/$exit
      -- CP-element group 57: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315__exit__
      -- CP-element group 57: 	 branch_block_stmt_1091/if_stmt_1316_dead_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1091/if_stmt_1316_eval_test/$entry
      -- CP-element group 57: 	 branch_block_stmt_1091/if_stmt_1316_eval_test/$exit
      -- CP-element group 57: 	 branch_block_stmt_1091/if_stmt_1316_eval_test/branch_req
      -- CP-element group 57: 	 branch_block_stmt_1091/R_exitcond1_1317_place
      -- CP-element group 57: 	 branch_block_stmt_1091/if_stmt_1316_if_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1091/if_stmt_1316_else_link/$entry
      -- 
    branch_req_3813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(57), ack => if_stmt_1316_branch_req_0); -- 
    sendOutput_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(12) & sendOutput_CP_3266_elements(56);
      gj_sendOutput_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  merge  transition  place  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	66 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1091/forx_xendx_xloopexit_forx_xend
      -- CP-element group 58: 	 branch_block_stmt_1091/merge_stmt_1322__exit__
      -- CP-element group 58: 	 branch_block_stmt_1091/if_stmt_1316_if_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1091/if_stmt_1316_if_link/if_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1091/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 58: 	 branch_block_stmt_1091/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1091/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1091/merge_stmt_1322_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1091/merge_stmt_1322_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1091/merge_stmt_1322_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1091/merge_stmt_1322_PhiAck/dummy
      -- CP-element group 58: 	 branch_block_stmt_1091/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1091/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_3818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1316_branch_ack_1, ack => sendOutput_CP_3266_elements(58)); -- 
    -- CP-element group 59:  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: 	62 
    -- CP-element group 59:  members (12) 
      -- CP-element group 59: 	 branch_block_stmt_1091/if_stmt_1316_else_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1091/if_stmt_1316_else_link/else_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1091/forx_xbody_forx_xbody
      -- CP-element group 59: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/$entry
      -- CP-element group 59: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/$entry
      -- CP-element group 59: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1316_branch_ack_0, ack => sendOutput_CP_3266_elements(59)); -- 
    rr_3866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(59), ack => type_cast_1194_inst_req_0); -- 
    cr_3871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(59), ack => type_cast_1194_inst_req_1); -- 
    -- CP-element group 60:  transition  output  delay-element  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	11 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	64 
    -- CP-element group 60:  members (5) 
      -- CP-element group 60: 	 branch_block_stmt_1091/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_1091/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1188/$exit
      -- CP-element group 60: 	 branch_block_stmt_1091/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/$exit
      -- CP-element group 60: 	 branch_block_stmt_1091/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1192_konst_delay_trans
      -- CP-element group 60: 	 branch_block_stmt_1091/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_req
      -- 
    phi_stmt_1188_req_3847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1188_req_3847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(60), ack => phi_stmt_1188_req_0); -- 
    -- Element group sendOutput_CP_3266_elements(60) is a control-delay.
    cp_element_60_delay: control_delay_element  generic map(name => " 60_delay", delay_value => 1)  port map(req => sendOutput_CP_3266_elements(11), ack => sendOutput_CP_3266_elements(60), clk => clk, reset =>reset);
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/SplitProtocol/Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/SplitProtocol/Sample/ra
      -- 
    ra_3867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1194_inst_ack_0, ack => sendOutput_CP_3266_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/SplitProtocol/Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/SplitProtocol/Update/ca
      -- 
    ca_3872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1194_inst_ack_1, ack => sendOutput_CP_3266_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/$exit
      -- CP-element group 63: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/$exit
      -- CP-element group 63: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/$exit
      -- CP-element group 63: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_sources/type_cast_1194/SplitProtocol/$exit
      -- CP-element group 63: 	 branch_block_stmt_1091/forx_xbody_forx_xbody_PhiReq/phi_stmt_1188/phi_stmt_1188_req
      -- 
    phi_stmt_1188_req_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1188_req_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(63), ack => phi_stmt_1188_req_1); -- 
    sendOutput_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(61) & sendOutput_CP_3266_elements(62);
      gj_sendOutput_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  merge  transition  place  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	60 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1091/merge_stmt_1187_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1091/merge_stmt_1187_PhiAck/$entry
      -- 
    sendOutput_CP_3266_elements(64) <= OrReduce(sendOutput_CP_3266_elements(60) & sendOutput_CP_3266_elements(63));
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	23 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	13 
    -- CP-element group 65: 	19 
    -- CP-element group 65: 	15 
    -- CP-element group 65: 	17 
    -- CP-element group 65: 	33 
    -- CP-element group 65: 	31 
    -- CP-element group 65: 	21 
    -- CP-element group 65: 	27 
    -- CP-element group 65: 	29 
    -- CP-element group 65: 	25 
    -- CP-element group 65:  members (53) 
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_scale_1/scale_rename_ack
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_resized_1
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_final_index_sum_regn_Update/req
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/word_access_complete/word_0/cr
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_final_index_sum_regn_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_scale_1/scale_rename_req
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_scale_1/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_scale_1/$exit
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1229_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_scaled_1
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_complete/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/addr_of_1201_complete/req
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1209_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_computed_1
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/word_access_complete/word_0/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_resize_1/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/merge_stmt_1187__exit__
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315__entry__
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_resize_1/$exit
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_Update/word_access_complete/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_resize_1/index_resize_req
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1249_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1219_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_index_resize_1/index_resize_ack
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/ptr_deref_1205_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_final_index_sum_regn_update_start
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1269_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1279_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_final_index_sum_regn_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1259_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/array_obj_ref_1200_final_index_sum_regn_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1091/assign_stmt_1202_to_assign_stmt_1315/type_cast_1239_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1091/merge_stmt_1187_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_1091/merge_stmt_1187_PhiAck/phi_stmt_1188_ack
      -- 
    phi_stmt_1188_ack_3878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1188_ack_0, ack => sendOutput_CP_3266_elements(65)); -- 
    req_3515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => array_obj_ref_1200_index_offset_req_1); -- 
    cr_3575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => ptr_deref_1205_load_0_req_1); -- 
    cr_3622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1229_inst_req_1); -- 
    cr_3594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1209_inst_req_1); -- 
    cr_3636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1239_inst_req_1); -- 
    req_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => addr_of_1201_final_reg_req_1); -- 
    cr_3692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1279_inst_req_1); -- 
    cr_3650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1249_inst_req_1); -- 
    cr_3608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1219_inst_req_1); -- 
    cr_3678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1269_inst_req_1); -- 
    req_3510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => array_obj_ref_1200_index_offset_req_0); -- 
    cr_3664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1259_inst_req_1); -- 
    -- CP-element group 66:  merge  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	9 
    -- CP-element group 66: 	58 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_1091/branch_block_stmt_1091__exit__
      -- CP-element group 66: 	 branch_block_stmt_1091/merge_stmt_1326__exit__
      -- CP-element group 66: 	 branch_block_stmt_1091/return__
      -- CP-element group 66: 	 branch_block_stmt_1091/merge_stmt_1324__exit__
      -- CP-element group 66: 	 branch_block_stmt_1091/$exit
      -- CP-element group 66: 	 $exit
      -- CP-element group 66: 	 branch_block_stmt_1091/merge_stmt_1324_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_1091/merge_stmt_1324_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_1091/merge_stmt_1324_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_1091/merge_stmt_1324_PhiAck/dummy
      -- CP-element group 66: 	 branch_block_stmt_1091/return___PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1091/return___PhiReq/$exit
      -- CP-element group 66: 	 branch_block_stmt_1091/merge_stmt_1326_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_1091/merge_stmt_1326_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_1091/merge_stmt_1326_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_1091/merge_stmt_1326_PhiAck/dummy
      -- 
    sendOutput_CP_3266_elements(66) <= OrReduce(sendOutput_CP_3266_elements(9) & sendOutput_CP_3266_elements(58));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_1199_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1199_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1200_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1200_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1200_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1200_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1200_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1200_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1202 : std_logic_vector(31 downto 0);
    signal cmp73_1143 : std_logic_vector(0 downto 0);
    signal conv17_1220 : std_logic_vector(7 downto 0);
    signal conv23_1230 : std_logic_vector(7 downto 0);
    signal conv29_1240 : std_logic_vector(7 downto 0);
    signal conv35_1250 : std_logic_vector(7 downto 0);
    signal conv41_1260 : std_logic_vector(7 downto 0);
    signal conv47_1270 : std_logic_vector(7 downto 0);
    signal conv53_1280 : std_logic_vector(7 downto 0);
    signal conv_1210 : std_logic_vector(7 downto 0);
    signal exitcond1_1315 : std_logic_vector(0 downto 0);
    signal iNsTr_0_1099 : std_logic_vector(31 downto 0);
    signal iNsTr_1_1111 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1123 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1172 : std_logic_vector(63 downto 0);
    signal indvar_1188 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1310 : std_logic_vector(63 downto 0);
    signal mul3_1137 : std_logic_vector(31 downto 0);
    signal mul_1132 : std_logic_vector(31 downto 0);
    signal ptr_deref_1102_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1102_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1102_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1102_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1102_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1114_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1114_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1114_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1114_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1114_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1126_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1126_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1126_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1126_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1126_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1205_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1205_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1205_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1205_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1205_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr14_1216 : std_logic_vector(63 downto 0);
    signal shr20_1226 : std_logic_vector(63 downto 0);
    signal shr26_1236 : std_logic_vector(63 downto 0);
    signal shr32_1246 : std_logic_vector(63 downto 0);
    signal shr38_1256 : std_logic_vector(63 downto 0);
    signal shr44_1266 : std_logic_vector(63 downto 0);
    signal shr50_1276 : std_logic_vector(63 downto 0);
    signal tmp1_1115 : std_logic_vector(31 downto 0);
    signal tmp2_1127 : std_logic_vector(31 downto 0);
    signal tmp77_1156 : std_logic_vector(31 downto 0);
    signal tmp77x_xop_1168 : std_logic_vector(31 downto 0);
    signal tmp78_1162 : std_logic_vector(0 downto 0);
    signal tmp81_1185 : std_logic_vector(63 downto 0);
    signal tmp9_1206 : std_logic_vector(63 downto 0);
    signal tmp_1103 : std_logic_vector(31 downto 0);
    signal type_cast_1141_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1154_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1160_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1166_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1176_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1183_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1192_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1194_wire : std_logic_vector(63 downto 0);
    signal type_cast_1214_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1224_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1234_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1244_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1254_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1264_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1274_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1308_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_1178 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1200_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1200_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1200_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1200_resized_base_address <= "00000000000000";
    iNsTr_0_1099 <= "00000000000000000000000000000010";
    iNsTr_1_1111 <= "00000000000000000000000000000011";
    iNsTr_2_1123 <= "00000000000000000000000000000100";
    ptr_deref_1102_word_offset_0 <= "0000000";
    ptr_deref_1114_word_offset_0 <= "0000000";
    ptr_deref_1126_word_offset_0 <= "0000000";
    ptr_deref_1205_word_offset_0 <= "00000000000000";
    type_cast_1141_wire_constant <= "00000000000000000000000000000011";
    type_cast_1154_wire_constant <= "00000000000000000000000000000010";
    type_cast_1160_wire_constant <= "00000000000000000000000000000001";
    type_cast_1166_wire_constant <= "11111111111111111111111111111111";
    type_cast_1176_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1183_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1192_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1214_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1224_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1234_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1244_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1254_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1264_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1274_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1308_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1188: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1192_wire_constant & type_cast_1194_wire;
      req <= phi_stmt_1188_req_0 & phi_stmt_1188_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1188",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1188_ack_0,
          idata => idata,
          odata => indvar_1188,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1188
    -- flow-through select operator MUX_1184_inst
    tmp81_1185 <= xx_xop_1178 when (tmp78_1162(0) /=  '0') else type_cast_1183_wire_constant;
    addr_of_1201_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1201_final_reg_req_0;
      addr_of_1201_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1201_final_reg_req_1;
      addr_of_1201_final_reg_ack_1<= rack(0);
      addr_of_1201_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1201_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1200_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1171_inst_req_0;
      type_cast_1171_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1171_inst_req_1;
      type_cast_1171_inst_ack_1<= rack(0);
      type_cast_1171_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1171_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp77x_xop_1168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_4_1172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1194_inst_req_0;
      type_cast_1194_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1194_inst_req_1;
      type_cast_1194_inst_ack_1<= rack(0);
      type_cast_1194_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1310,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1194_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1209_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1209_inst_req_0;
      type_cast_1209_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1209_inst_req_1;
      type_cast_1209_inst_ack_1<= rack(0);
      type_cast_1209_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1209_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp9_1206,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1219_inst_req_0;
      type_cast_1219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1219_inst_req_1;
      type_cast_1219_inst_ack_1<= rack(0);
      type_cast_1219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr14_1216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1229_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1229_inst_req_0;
      type_cast_1229_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1229_inst_req_1;
      type_cast_1229_inst_ack_1<= rack(0);
      type_cast_1229_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1229_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr20_1226,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_1230,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1239_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1239_inst_req_0;
      type_cast_1239_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1239_inst_req_1;
      type_cast_1239_inst_ack_1<= rack(0);
      type_cast_1239_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1239_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr26_1236,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1240,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1249_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1249_inst_req_0;
      type_cast_1249_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1249_inst_req_1;
      type_cast_1249_inst_ack_1<= rack(0);
      type_cast_1249_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1249_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr32_1246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_1250,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1259_inst_req_0;
      type_cast_1259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1259_inst_req_1;
      type_cast_1259_inst_ack_1<= rack(0);
      type_cast_1259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr38_1256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_1260,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1269_inst_req_0;
      type_cast_1269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1269_inst_req_1;
      type_cast_1269_inst_ack_1<= rack(0);
      type_cast_1269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr44_1266,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_1270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1279_inst_req_0;
      type_cast_1279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1279_inst_req_1;
      type_cast_1279_inst_ack_1<= rack(0);
      type_cast_1279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr50_1276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_1280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1200_index_1_rename
    process(R_indvar_1199_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1199_resized;
      ov(13 downto 0) := iv;
      R_indvar_1199_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1200_index_1_resize
    process(indvar_1188) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1188;
      ov := iv(13 downto 0);
      R_indvar_1199_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1200_root_address_inst
    process(array_obj_ref_1200_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1200_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1200_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1102_addr_0
    process(ptr_deref_1102_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1102_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1102_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1102_base_resize
    process(iNsTr_0_1099) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_1099;
      ov := iv(6 downto 0);
      ptr_deref_1102_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1102_gather_scatter
    process(ptr_deref_1102_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1102_data_0;
      ov(31 downto 0) := iv;
      tmp_1103 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1102_root_address_inst
    process(ptr_deref_1102_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1102_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1102_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1114_addr_0
    process(ptr_deref_1114_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1114_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1114_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1114_base_resize
    process(iNsTr_1_1111) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_1111;
      ov := iv(6 downto 0);
      ptr_deref_1114_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1114_gather_scatter
    process(ptr_deref_1114_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1114_data_0;
      ov(31 downto 0) := iv;
      tmp1_1115 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1114_root_address_inst
    process(ptr_deref_1114_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1114_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1114_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1126_addr_0
    process(ptr_deref_1126_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1126_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1126_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1126_base_resize
    process(iNsTr_2_1123) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1123;
      ov := iv(6 downto 0);
      ptr_deref_1126_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1126_gather_scatter
    process(ptr_deref_1126_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1126_data_0;
      ov(31 downto 0) := iv;
      tmp2_1127 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1126_root_address_inst
    process(ptr_deref_1126_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1126_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1126_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1205_addr_0
    process(ptr_deref_1205_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1205_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1205_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1205_base_resize
    process(arrayidx_1202) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1202;
      ov := iv(13 downto 0);
      ptr_deref_1205_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1205_gather_scatter
    process(ptr_deref_1205_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1205_data_0;
      ov(63 downto 0) := iv;
      tmp9_1206 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1205_root_address_inst
    process(ptr_deref_1205_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1205_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1205_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1144_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp73_1143;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1144_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1144_branch_req_0,
          ack0 => if_stmt_1144_branch_ack_0,
          ack1 => if_stmt_1144_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1316_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1315;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1316_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1316_branch_req_0,
          ack0 => if_stmt_1316_branch_ack_0,
          ack1 => if_stmt_1316_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1167_inst
    process(tmp77_1156) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp77_1156, type_cast_1166_wire_constant, tmp_var);
      tmp77x_xop_1168 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1177_inst
    process(iNsTr_4_1172) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_4_1172, type_cast_1176_wire_constant, tmp_var);
      xx_xop_1178 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1309_inst
    process(indvar_1188) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1188, type_cast_1308_wire_constant, tmp_var);
      indvarx_xnext_1310 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1314_inst
    process(indvarx_xnext_1310, tmp81_1185) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1310, tmp81_1185, tmp_var);
      exitcond1_1315 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1155_inst
    process(mul3_1137) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul3_1137, type_cast_1154_wire_constant, tmp_var);
      tmp77_1156 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1215_inst
    process(tmp9_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1206, type_cast_1214_wire_constant, tmp_var);
      shr14_1216 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1225_inst
    process(tmp9_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1206, type_cast_1224_wire_constant, tmp_var);
      shr20_1226 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1235_inst
    process(tmp9_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1206, type_cast_1234_wire_constant, tmp_var);
      shr26_1236 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1245_inst
    process(tmp9_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1206, type_cast_1244_wire_constant, tmp_var);
      shr32_1246 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1255_inst
    process(tmp9_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1206, type_cast_1254_wire_constant, tmp_var);
      shr38_1256 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1265_inst
    process(tmp9_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1206, type_cast_1264_wire_constant, tmp_var);
      shr44_1266 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1275_inst
    process(tmp9_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1206, type_cast_1274_wire_constant, tmp_var);
      shr50_1276 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1131_inst
    process(tmp1_1115, tmp_1103) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_1115, tmp_1103, tmp_var);
      mul_1132 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1136_inst
    process(mul_1132, tmp2_1127) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1132, tmp2_1127, tmp_var);
      mul3_1137 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1142_inst
    process(mul3_1137) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul3_1137, type_cast_1141_wire_constant, tmp_var);
      cmp73_1143 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1161_inst
    process(tmp77_1156) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp77_1156, type_cast_1160_wire_constant, tmp_var);
      tmp78_1162 <= tmp_var; --
    end process;
    -- shared split operator group (16) : array_obj_ref_1200_index_offset 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1199_scaled;
      array_obj_ref_1200_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1200_index_offset_req_0;
      array_obj_ref_1200_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1200_index_offset_req_1;
      array_obj_ref_1200_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared load operator group (0) : ptr_deref_1102_load_0 ptr_deref_1114_load_0 ptr_deref_1126_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1102_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1114_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1126_load_0_req_0;
      ptr_deref_1102_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1114_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1126_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1102_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1114_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1126_load_0_req_1;
      ptr_deref_1102_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1114_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1126_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1102_word_address_0 & ptr_deref_1114_word_address_0 & ptr_deref_1126_word_address_0;
      ptr_deref_1102_data_0 <= data_out(95 downto 64);
      ptr_deref_1114_data_0 <= data_out(63 downto 32);
      ptr_deref_1126_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1205_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1205_load_0_req_0;
      ptr_deref_1205_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1205_load_0_req_1;
      ptr_deref_1205_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1205_word_address_0;
      ptr_deref_1205_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(13 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(63 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_1296_inst WPIPE_ConvTranspose_output_pipe_1290_inst WPIPE_ConvTranspose_output_pipe_1299_inst WPIPE_ConvTranspose_output_pipe_1293_inst WPIPE_ConvTranspose_output_pipe_1287_inst WPIPE_ConvTranspose_output_pipe_1284_inst WPIPE_ConvTranspose_output_pipe_1281_inst WPIPE_ConvTranspose_output_pipe_1302_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1296_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1290_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1299_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1293_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1287_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1284_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1281_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1302_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1296_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1290_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1299_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1293_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1287_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1284_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1281_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1302_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv23_1230 & conv35_1250 & conv17_1220 & conv29_1240 & conv41_1260 & conv47_1270 & conv53_1280 & conv_1210;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_0_start: Boolean;
  signal testConfigure_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_468_load_0_ack_1 : boolean;
  signal ptr_deref_468_load_0_ack_0 : boolean;
  signal type_cast_487_inst_ack_1 : boolean;
  signal ptr_deref_468_load_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_ack_1 : boolean;
  signal type_cast_861_inst_req_1 : boolean;
  signal if_stmt_501_branch_ack_1 : boolean;
  signal if_stmt_501_branch_ack_0 : boolean;
  signal if_stmt_501_branch_req_0 : boolean;
  signal if_stmt_937_branch_ack_1 : boolean;
  signal type_cast_861_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_857_inst_req_0 : boolean;
  signal ptr_deref_369_store_0_ack_0 : boolean;
  signal ptr_deref_369_store_0_req_0 : boolean;
  signal ptr_deref_382_load_0_req_0 : boolean;
  signal type_cast_358_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_875_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 : boolean;
  signal ptr_deref_456_load_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 : boolean;
  signal ptr_deref_468_load_0_req_0 : boolean;
  signal ptr_deref_432_load_0_req_0 : boolean;
  signal type_cast_39_inst_req_0 : boolean;
  signal type_cast_39_inst_ack_0 : boolean;
  signal type_cast_39_inst_req_1 : boolean;
  signal type_cast_39_inst_ack_1 : boolean;
  signal ptr_deref_456_load_0_req_1 : boolean;
  signal ptr_deref_444_load_0_ack_1 : boolean;
  signal ptr_deref_48_store_0_req_0 : boolean;
  signal ptr_deref_48_store_0_ack_0 : boolean;
  signal ptr_deref_48_store_0_req_1 : boolean;
  signal ptr_deref_48_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 : boolean;
  signal if_stmt_998_branch_req_0 : boolean;
  signal type_cast_63_inst_req_0 : boolean;
  signal type_cast_897_inst_ack_0 : boolean;
  signal type_cast_63_inst_ack_0 : boolean;
  signal ptr_deref_444_load_0_req_1 : boolean;
  signal type_cast_63_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_1 : boolean;
  signal type_cast_487_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_857_inst_ack_0 : boolean;
  signal if_stmt_65_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_857_inst_ack_1 : boolean;
  signal if_stmt_65_branch_ack_1 : boolean;
  signal ptr_deref_406_load_0_ack_1 : boolean;
  signal if_stmt_65_branch_ack_0 : boolean;
  signal ptr_deref_406_load_0_req_1 : boolean;
  signal type_cast_96_inst_req_0 : boolean;
  signal type_cast_96_inst_ack_0 : boolean;
  signal type_cast_96_inst_req_1 : boolean;
  signal type_cast_96_inst_ack_1 : boolean;
  signal type_cast_487_inst_req_0 : boolean;
  signal ptr_deref_432_load_0_ack_1 : boolean;
  signal ptr_deref_432_load_0_req_1 : boolean;
  signal array_obj_ref_102_index_offset_req_0 : boolean;
  signal array_obj_ref_102_index_offset_ack_0 : boolean;
  signal array_obj_ref_102_index_offset_req_1 : boolean;
  signal array_obj_ref_102_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_857_inst_req_1 : boolean;
  signal addr_of_103_final_reg_req_0 : boolean;
  signal addr_of_103_final_reg_ack_0 : boolean;
  signal addr_of_103_final_reg_req_1 : boolean;
  signal addr_of_103_final_reg_ack_1 : boolean;
  signal ptr_deref_432_load_0_ack_0 : boolean;
  signal ptr_deref_456_load_0_ack_0 : boolean;
  signal type_cast_897_inst_req_1 : boolean;
  signal type_cast_1025_inst_req_0 : boolean;
  signal ptr_deref_456_load_0_req_0 : boolean;
  signal ptr_deref_106_store_0_req_0 : boolean;
  signal ptr_deref_106_store_0_ack_0 : boolean;
  signal ptr_deref_106_store_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_875_inst_req_0 : boolean;
  signal ptr_deref_106_store_0_ack_1 : boolean;
  signal type_cast_420_inst_ack_1 : boolean;
  signal addr_of_275_final_reg_req_0 : boolean;
  signal addr_of_275_final_reg_ack_0 : boolean;
  signal addr_of_275_final_reg_req_1 : boolean;
  signal addr_of_275_final_reg_ack_1 : boolean;
  signal ptr_deref_369_store_0_ack_1 : boolean;
  signal ptr_deref_394_load_0_ack_0 : boolean;
  signal type_cast_420_inst_req_1 : boolean;
  signal ptr_deref_123_load_0_req_0 : boolean;
  signal ptr_deref_123_load_0_ack_0 : boolean;
  signal ptr_deref_123_load_0_req_1 : boolean;
  signal ptr_deref_123_load_0_ack_1 : boolean;
  signal type_cast_358_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_131_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_131_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_131_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_131_inst_ack_1 : boolean;
  signal ptr_deref_444_load_0_ack_0 : boolean;
  signal type_cast_135_inst_req_0 : boolean;
  signal type_cast_135_inst_ack_0 : boolean;
  signal type_cast_135_inst_req_1 : boolean;
  signal type_cast_135_inst_ack_1 : boolean;
  signal if_stmt_937_branch_ack_0 : boolean;
  signal type_cast_1025_inst_ack_0 : boolean;
  signal ptr_deref_444_load_0_req_0 : boolean;
  signal if_stmt_137_branch_req_0 : boolean;
  signal type_cast_358_inst_req_1 : boolean;
  signal if_stmt_137_branch_ack_1 : boolean;
  signal if_stmt_137_branch_ack_0 : boolean;
  signal type_cast_420_inst_ack_0 : boolean;
  signal type_cast_915_inst_req_0 : boolean;
  signal type_cast_420_inst_req_0 : boolean;
  signal ptr_deref_165_store_0_req_0 : boolean;
  signal ptr_deref_165_store_0_ack_0 : boolean;
  signal ptr_deref_165_store_0_req_1 : boolean;
  signal ptr_deref_165_store_0_ack_1 : boolean;
  signal ptr_deref_406_load_0_ack_0 : boolean;
  signal if_stmt_174_branch_req_0 : boolean;
  signal if_stmt_174_branch_ack_1 : boolean;
  signal ptr_deref_406_load_0_req_0 : boolean;
  signal if_stmt_174_branch_ack_0 : boolean;
  signal ptr_deref_382_load_0_ack_1 : boolean;
  signal type_cast_199_inst_req_0 : boolean;
  signal type_cast_199_inst_ack_0 : boolean;
  signal type_cast_199_inst_req_1 : boolean;
  signal type_cast_199_inst_ack_1 : boolean;
  signal array_obj_ref_205_index_offset_req_0 : boolean;
  signal array_obj_ref_205_index_offset_ack_0 : boolean;
  signal array_obj_ref_205_index_offset_req_1 : boolean;
  signal array_obj_ref_205_index_offset_ack_1 : boolean;
  signal addr_of_206_final_reg_req_0 : boolean;
  signal type_cast_915_inst_ack_0 : boolean;
  signal addr_of_206_final_reg_ack_0 : boolean;
  signal addr_of_206_final_reg_req_1 : boolean;
  signal addr_of_206_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_209_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_209_inst_ack_0 : boolean;
  signal ptr_deref_382_load_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_209_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_209_inst_ack_1 : boolean;
  signal type_cast_213_inst_req_0 : boolean;
  signal type_cast_213_inst_ack_0 : boolean;
  signal type_cast_213_inst_req_1 : boolean;
  signal type_cast_213_inst_ack_1 : boolean;
  signal ptr_deref_216_store_0_req_0 : boolean;
  signal ptr_deref_216_store_0_ack_0 : boolean;
  signal ptr_deref_216_store_0_req_1 : boolean;
  signal ptr_deref_216_store_0_ack_1 : boolean;
  signal type_cast_897_inst_req_0 : boolean;
  signal ptr_deref_233_load_0_req_0 : boolean;
  signal ptr_deref_233_load_0_ack_0 : boolean;
  signal ptr_deref_382_load_0_ack_0 : boolean;
  signal ptr_deref_233_load_0_req_1 : boolean;
  signal ptr_deref_233_load_0_ack_1 : boolean;
  signal type_cast_487_inst_req_1 : boolean;
  signal type_cast_897_inst_ack_1 : boolean;
  signal if_stmt_240_branch_req_0 : boolean;
  signal if_stmt_240_branch_ack_1 : boolean;
  signal type_cast_358_inst_req_0 : boolean;
  signal if_stmt_240_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_250_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_250_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_250_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_250_inst_ack_1 : boolean;
  signal type_cast_254_inst_req_0 : boolean;
  signal type_cast_254_inst_ack_0 : boolean;
  signal type_cast_254_inst_req_1 : boolean;
  signal type_cast_254_inst_ack_1 : boolean;
  signal type_cast_1025_inst_req_1 : boolean;
  signal ptr_deref_394_load_0_ack_1 : boolean;
  signal ptr_deref_394_load_0_req_1 : boolean;
  signal ptr_deref_369_store_0_req_1 : boolean;
  signal ptr_deref_394_load_0_req_0 : boolean;
  signal ptr_deref_278_store_0_req_0 : boolean;
  signal ptr_deref_278_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_875_inst_ack_0 : boolean;
  signal ptr_deref_278_store_0_req_1 : boolean;
  signal ptr_deref_278_store_0_ack_1 : boolean;
  signal type_cast_1025_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_req_0 : boolean;
  signal ptr_deref_980_load_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_ack_1 : boolean;
  signal type_cast_286_inst_req_0 : boolean;
  signal type_cast_286_inst_ack_0 : boolean;
  signal type_cast_286_inst_req_1 : boolean;
  signal type_cast_286_inst_ack_1 : boolean;
  signal if_stmt_998_branch_ack_1 : boolean;
  signal if_stmt_300_branch_req_0 : boolean;
  signal if_stmt_300_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_875_inst_req_1 : boolean;
  signal if_stmt_300_branch_ack_0 : boolean;
  signal ptr_deref_980_load_0_ack_0 : boolean;
  signal addr_of_1055_final_reg_req_0 : boolean;
  signal STORE_padding_312_store_0_req_0 : boolean;
  signal STORE_padding_312_store_0_ack_0 : boolean;
  signal type_cast_915_inst_req_1 : boolean;
  signal STORE_padding_312_store_0_req_1 : boolean;
  signal STORE_padding_312_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_911_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_911_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 : boolean;
  signal ptr_deref_956_load_0_req_0 : boolean;
  signal addr_of_1055_final_reg_ack_0 : boolean;
  signal ptr_deref_956_load_0_ack_0 : boolean;
  signal type_cast_915_inst_ack_1 : boolean;
  signal type_cast_320_inst_req_0 : boolean;
  signal type_cast_320_inst_ack_0 : boolean;
  signal type_cast_320_inst_req_1 : boolean;
  signal type_cast_320_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_911_inst_req_1 : boolean;
  signal ptr_deref_331_store_0_req_0 : boolean;
  signal ptr_deref_331_store_0_ack_0 : boolean;
  signal ptr_deref_331_store_0_req_1 : boolean;
  signal ptr_deref_331_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_ack_1 : boolean;
  signal type_cast_339_inst_req_0 : boolean;
  signal type_cast_339_inst_ack_0 : boolean;
  signal type_cast_339_inst_req_1 : boolean;
  signal type_cast_339_inst_ack_1 : boolean;
  signal ptr_deref_350_store_0_req_0 : boolean;
  signal ptr_deref_350_store_0_ack_0 : boolean;
  signal ptr_deref_350_store_0_req_1 : boolean;
  signal ptr_deref_350_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_req_1 : boolean;
  signal type_cast_843_inst_ack_1 : boolean;
  signal if_stmt_522_branch_req_0 : boolean;
  signal type_cast_861_inst_ack_0 : boolean;
  signal if_stmt_522_branch_ack_1 : boolean;
  signal if_stmt_522_branch_ack_0 : boolean;
  signal type_cast_541_inst_req_0 : boolean;
  signal type_cast_541_inst_ack_0 : boolean;
  signal type_cast_541_inst_req_1 : boolean;
  signal type_cast_541_inst_ack_1 : boolean;
  signal if_stmt_937_branch_req_0 : boolean;
  signal type_cast_861_inst_req_0 : boolean;
  signal array_obj_ref_576_index_offset_req_0 : boolean;
  signal array_obj_ref_576_index_offset_ack_0 : boolean;
  signal array_obj_ref_576_index_offset_req_1 : boolean;
  signal array_obj_ref_576_index_offset_ack_1 : boolean;
  signal addr_of_577_final_reg_req_0 : boolean;
  signal addr_of_577_final_reg_ack_0 : boolean;
  signal addr_of_577_final_reg_req_1 : boolean;
  signal addr_of_577_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_ack_0 : boolean;
  signal ptr_deref_923_store_0_ack_1 : boolean;
  signal ptr_deref_923_store_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_580_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_580_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_580_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_580_inst_ack_1 : boolean;
  signal type_cast_584_inst_req_0 : boolean;
  signal type_cast_584_inst_ack_0 : boolean;
  signal type_cast_584_inst_req_1 : boolean;
  signal type_cast_584_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_ack_1 : boolean;
  signal array_obj_ref_1054_index_offset_ack_1 : boolean;
  signal type_cast_597_inst_req_0 : boolean;
  signal type_cast_597_inst_ack_0 : boolean;
  signal type_cast_597_inst_req_1 : boolean;
  signal type_cast_597_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_ack_1 : boolean;
  signal ptr_deref_923_store_0_ack_0 : boolean;
  signal array_obj_ref_1054_index_offset_req_1 : boolean;
  signal type_cast_615_inst_req_0 : boolean;
  signal type_cast_615_inst_ack_0 : boolean;
  signal type_cast_615_inst_req_1 : boolean;
  signal type_cast_615_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_629_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_629_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_629_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_629_inst_ack_1 : boolean;
  signal ptr_deref_923_store_0_req_0 : boolean;
  signal type_cast_633_inst_req_0 : boolean;
  signal type_cast_633_inst_ack_0 : boolean;
  signal type_cast_633_inst_req_1 : boolean;
  signal type_cast_633_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_647_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_647_inst_ack_0 : boolean;
  signal type_cast_879_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_647_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_647_inst_ack_1 : boolean;
  signal type_cast_651_inst_req_0 : boolean;
  signal type_cast_651_inst_ack_0 : boolean;
  signal type_cast_651_inst_req_1 : boolean;
  signal type_cast_651_inst_ack_1 : boolean;
  signal addr_of_1055_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_665_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_665_inst_ack_0 : boolean;
  signal type_cast_879_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_665_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_665_inst_ack_1 : boolean;
  signal array_obj_ref_1054_index_offset_ack_0 : boolean;
  signal type_cast_669_inst_req_0 : boolean;
  signal type_cast_669_inst_ack_0 : boolean;
  signal type_cast_669_inst_req_1 : boolean;
  signal type_cast_669_inst_ack_1 : boolean;
  signal addr_of_1055_final_reg_req_1 : boolean;
  signal if_stmt_998_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_683_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_683_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_683_inst_req_1 : boolean;
  signal ptr_deref_968_load_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_683_inst_ack_1 : boolean;
  signal array_obj_ref_1054_index_offset_req_0 : boolean;
  signal type_cast_687_inst_req_0 : boolean;
  signal ptr_deref_968_load_0_req_1 : boolean;
  signal type_cast_687_inst_ack_0 : boolean;
  signal type_cast_687_inst_req_1 : boolean;
  signal type_cast_687_inst_ack_1 : boolean;
  signal type_cast_879_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_701_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_701_inst_ack_0 : boolean;
  signal type_cast_879_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_701_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_701_inst_ack_1 : boolean;
  signal type_cast_705_inst_req_0 : boolean;
  signal type_cast_705_inst_ack_0 : boolean;
  signal type_cast_705_inst_req_1 : boolean;
  signal type_cast_705_inst_ack_1 : boolean;
  signal ptr_deref_1058_store_0_req_0 : boolean;
  signal ptr_deref_980_load_0_ack_1 : boolean;
  signal ptr_deref_980_load_0_req_1 : boolean;
  signal ptr_deref_968_load_0_ack_0 : boolean;
  signal ptr_deref_968_load_0_req_0 : boolean;
  signal ptr_deref_713_store_0_req_0 : boolean;
  signal ptr_deref_713_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_911_inst_ack_1 : boolean;
  signal ptr_deref_713_store_0_req_1 : boolean;
  signal ptr_deref_713_store_0_ack_1 : boolean;
  signal type_cast_843_inst_req_1 : boolean;
  signal ptr_deref_956_load_0_ack_1 : boolean;
  signal if_stmt_727_branch_req_0 : boolean;
  signal ptr_deref_956_load_0_req_1 : boolean;
  signal if_stmt_727_branch_ack_1 : boolean;
  signal if_stmt_727_branch_ack_0 : boolean;
  signal type_cast_751_inst_req_0 : boolean;
  signal type_cast_751_inst_ack_0 : boolean;
  signal type_cast_751_inst_req_1 : boolean;
  signal type_cast_751_inst_ack_1 : boolean;
  signal array_obj_ref_786_index_offset_req_0 : boolean;
  signal array_obj_ref_786_index_offset_ack_0 : boolean;
  signal array_obj_ref_786_index_offset_req_1 : boolean;
  signal array_obj_ref_786_index_offset_ack_1 : boolean;
  signal addr_of_787_final_reg_req_0 : boolean;
  signal addr_of_787_final_reg_ack_0 : boolean;
  signal addr_of_787_final_reg_req_1 : boolean;
  signal addr_of_787_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_790_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_790_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_790_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_790_inst_ack_1 : boolean;
  signal type_cast_794_inst_req_0 : boolean;
  signal type_cast_794_inst_ack_0 : boolean;
  signal type_cast_794_inst_req_1 : boolean;
  signal type_cast_794_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_803_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_803_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_803_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_803_inst_ack_1 : boolean;
  signal type_cast_807_inst_req_0 : boolean;
  signal type_cast_807_inst_ack_0 : boolean;
  signal type_cast_807_inst_req_1 : boolean;
  signal type_cast_807_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_821_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_821_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_821_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_821_inst_ack_1 : boolean;
  signal type_cast_825_inst_req_0 : boolean;
  signal type_cast_825_inst_ack_0 : boolean;
  signal type_cast_825_inst_req_1 : boolean;
  signal type_cast_825_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_839_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_839_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_839_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_839_inst_ack_1 : boolean;
  signal type_cast_843_inst_req_0 : boolean;
  signal type_cast_843_inst_ack_0 : boolean;
  signal ptr_deref_1058_store_0_ack_0 : boolean;
  signal ptr_deref_1058_store_0_req_1 : boolean;
  signal ptr_deref_1058_store_0_ack_1 : boolean;
  signal if_stmt_1073_branch_req_0 : boolean;
  signal if_stmt_1073_branch_ack_1 : boolean;
  signal if_stmt_1073_branch_ack_0 : boolean;
  signal type_cast_1084_inst_req_0 : boolean;
  signal type_cast_1084_inst_ack_0 : boolean;
  signal type_cast_1084_inst_req_1 : boolean;
  signal type_cast_1084_inst_ack_1 : boolean;
  signal type_cast_77_inst_req_0 : boolean;
  signal type_cast_77_inst_ack_0 : boolean;
  signal type_cast_77_inst_req_1 : boolean;
  signal type_cast_77_inst_ack_1 : boolean;
  signal phi_stmt_74_req_0 : boolean;
  signal type_cast_84_inst_req_0 : boolean;
  signal type_cast_84_inst_ack_0 : boolean;
  signal type_cast_84_inst_req_1 : boolean;
  signal type_cast_84_inst_ack_1 : boolean;
  signal phi_stmt_81_req_0 : boolean;
  signal phi_stmt_74_req_1 : boolean;
  signal type_cast_86_inst_req_0 : boolean;
  signal type_cast_86_inst_ack_0 : boolean;
  signal type_cast_86_inst_req_1 : boolean;
  signal type_cast_86_inst_ack_1 : boolean;
  signal phi_stmt_81_req_1 : boolean;
  signal phi_stmt_74_ack_0 : boolean;
  signal phi_stmt_81_ack_0 : boolean;
  signal type_cast_147_inst_req_0 : boolean;
  signal type_cast_147_inst_ack_0 : boolean;
  signal type_cast_147_inst_req_1 : boolean;
  signal type_cast_147_inst_ack_1 : boolean;
  signal phi_stmt_144_req_0 : boolean;
  signal phi_stmt_144_ack_0 : boolean;
  signal type_cast_154_inst_req_0 : boolean;
  signal type_cast_154_inst_ack_0 : boolean;
  signal type_cast_154_inst_req_1 : boolean;
  signal type_cast_154_inst_ack_1 : boolean;
  signal phi_stmt_151_req_0 : boolean;
  signal type_cast_156_inst_req_0 : boolean;
  signal type_cast_156_inst_ack_0 : boolean;
  signal type_cast_156_inst_req_1 : boolean;
  signal type_cast_156_inst_ack_1 : boolean;
  signal phi_stmt_151_req_1 : boolean;
  signal phi_stmt_151_ack_0 : boolean;
  signal type_cast_186_inst_req_0 : boolean;
  signal type_cast_186_inst_ack_0 : boolean;
  signal type_cast_186_inst_req_1 : boolean;
  signal type_cast_186_inst_ack_1 : boolean;
  signal phi_stmt_183_req_0 : boolean;
  signal phi_stmt_183_req_1 : boolean;
  signal phi_stmt_183_ack_0 : boolean;
  signal phi_stmt_258_req_0 : boolean;
  signal type_cast_268_inst_req_0 : boolean;
  signal type_cast_268_inst_ack_0 : boolean;
  signal type_cast_268_inst_req_1 : boolean;
  signal type_cast_268_inst_ack_1 : boolean;
  signal phi_stmt_265_req_0 : boolean;
  signal type_cast_264_inst_req_0 : boolean;
  signal type_cast_264_inst_ack_0 : boolean;
  signal type_cast_264_inst_req_1 : boolean;
  signal type_cast_264_inst_ack_1 : boolean;
  signal phi_stmt_258_req_1 : boolean;
  signal type_cast_270_inst_req_0 : boolean;
  signal type_cast_270_inst_ack_0 : boolean;
  signal type_cast_270_inst_req_1 : boolean;
  signal type_cast_270_inst_ack_1 : boolean;
  signal phi_stmt_265_req_1 : boolean;
  signal phi_stmt_258_ack_0 : boolean;
  signal phi_stmt_265_ack_0 : boolean;
  signal type_cast_310_inst_req_0 : boolean;
  signal type_cast_310_inst_ack_0 : boolean;
  signal type_cast_310_inst_req_1 : boolean;
  signal type_cast_310_inst_ack_1 : boolean;
  signal phi_stmt_307_req_0 : boolean;
  signal phi_stmt_307_ack_0 : boolean;
  signal phi_stmt_564_req_0 : boolean;
  signal type_cast_570_inst_req_0 : boolean;
  signal type_cast_570_inst_ack_0 : boolean;
  signal type_cast_570_inst_req_1 : boolean;
  signal type_cast_570_inst_ack_1 : boolean;
  signal phi_stmt_564_req_1 : boolean;
  signal phi_stmt_564_ack_0 : boolean;
  signal phi_stmt_774_req_0 : boolean;
  signal type_cast_780_inst_req_0 : boolean;
  signal type_cast_780_inst_ack_0 : boolean;
  signal type_cast_780_inst_req_1 : boolean;
  signal type_cast_780_inst_ack_1 : boolean;
  signal phi_stmt_774_req_1 : boolean;
  signal phi_stmt_774_ack_0 : boolean;
  signal phi_stmt_1042_req_0 : boolean;
  signal type_cast_1048_inst_req_0 : boolean;
  signal type_cast_1048_inst_ack_0 : boolean;
  signal type_cast_1048_inst_req_1 : boolean;
  signal type_cast_1048_inst_ack_1 : boolean;
  signal phi_stmt_1042_req_1 : boolean;
  signal phi_stmt_1042_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_0: Block -- control-path 
    signal testConfigure_CP_0_elements: BooleanArray(310 downto 0);
    -- 
  begin -- 
    testConfigure_CP_0_elements(0) <= testConfigure_CP_0_start;
    testConfigure_CP_0_symbol <= testConfigure_CP_0_elements(233);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (35) 
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_33/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/branch_block_stmt_33__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_Update/cr
      -- 
    rr_118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_0); -- 
    cr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_39_inst_req_1); -- 
    cr_187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => ptr_deref_48_store_0_req_1); -- 
    cr_215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_63_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_update_start_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_Update/cr
      -- 
    ra_119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_0, ack => testConfigure_CP_0_elements(1)); -- 
    cr_123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(1), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_35_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_Sample/rr
      -- 
    ca_124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_1, ack => testConfigure_CP_0_elements(2)); -- 
    rr_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => type_cast_39_inst_req_0); -- 
    rr_196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_Sample/ra
      -- 
    ra_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_39_inst_ack_0, ack => testConfigure_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_39_Update/ca
      -- 
    ca_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_39_inst_ack_1, ack => testConfigure_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/ptr_deref_48_Split/$entry
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/ptr_deref_48_Split/$exit
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/ptr_deref_48_Split/split_req
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/ptr_deref_48_Split/split_ack
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/word_access_start/$entry
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/word_access_start/word_0/rr
      -- 
    rr_176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(5), ack => ptr_deref_48_store_0_req_0); -- 
    testConfigure_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(0) & testConfigure_CP_0_elements(4);
      gj_testConfigure_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Sample/word_access_start/word_0/ra
      -- 
    ra_177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_48_store_0_ack_0, ack => testConfigure_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/ptr_deref_48_Update/word_access_complete/word_0/ca
      -- 
    ca_188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_48_store_0_ack_1, ack => testConfigure_CP_0_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_update_start_
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_Update/cr
      -- 
    ra_197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_0, ack => testConfigure_CP_0_elements(8)); -- 
    cr_201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(8), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/RPIPE_ConvTranspose_input_pipe_59_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_Sample/rr
      -- 
    ca_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_1, ack => testConfigure_CP_0_elements(9)); -- 
    rr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(9), ack => type_cast_63_inst_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_Sample/ra
      -- 
    ra_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_0, ack => testConfigure_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/type_cast_63_Update/ca
      -- 
    ca_216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_1, ack => testConfigure_CP_0_elements(11)); -- 
    -- CP-element group 12:  branch  join  transition  place  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (10) 
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64__exit__
      -- CP-element group 12: 	 branch_block_stmt_33/if_stmt_65__entry__
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_64/$exit
      -- CP-element group 12: 	 branch_block_stmt_33/if_stmt_65_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_33/if_stmt_65_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_33/if_stmt_65_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_33/if_stmt_65_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_33/R_cmp227_66_place
      -- CP-element group 12: 	 branch_block_stmt_33/if_stmt_65_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_33/if_stmt_65_else_link/$entry
      -- 
    branch_req_224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(12), ack => if_stmt_65_branch_req_0); -- 
    testConfigure_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(7) & testConfigure_CP_0_elements(11);
      gj_testConfigure_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	254 
    -- CP-element group 13: 	255 
    -- CP-element group 13:  members (12) 
      -- CP-element group 13: 	 branch_block_stmt_33/if_stmt_65_if_link/$exit
      -- CP-element group 13: 	 branch_block_stmt_33/if_stmt_65_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_33/entry_forx_xend
      -- CP-element group 13: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/SplitProtocol/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/SplitProtocol/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/SplitProtocol/Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/SplitProtocol/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/SplitProtocol/Update/cr
      -- 
    if_choice_transition_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_65_branch_ack_1, ack => testConfigure_CP_0_elements(13)); -- 
    rr_2787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_154_inst_req_0); -- 
    cr_2792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_154_inst_req_1); -- 
    -- CP-element group 14:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	241 
    -- CP-element group 14: 	242 
    -- CP-element group 14: 	243 
    -- CP-element group 14:  members (22) 
      -- CP-element group 14: 	 branch_block_stmt_33/merge_stmt_71__exit__
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody
      -- CP-element group 14: 	 branch_block_stmt_33/if_stmt_65_else_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_33/if_stmt_65_else_link/else_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_33/entry_forx_xbodyx_xpreheader
      -- CP-element group 14: 	 branch_block_stmt_33/entry_forx_xbodyx_xpreheader_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/entry_forx_xbodyx_xpreheader_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_33/merge_stmt_71_PhiReqMerge
      -- CP-element group 14: 	 branch_block_stmt_33/merge_stmt_71_PhiAck/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/merge_stmt_71_PhiAck/$exit
      -- CP-element group 14: 	 branch_block_stmt_33/merge_stmt_71_PhiAck/dummy
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_74/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/SplitProtocol/Update/cr
      -- 
    else_choice_transition_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_65_branch_ack_0, ack => testConfigure_CP_0_elements(14)); -- 
    rr_2720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_86_inst_req_0); -- 
    cr_2725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_86_inst_req_1); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	249 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_Sample/ra
      -- 
    ra_247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_96_inst_ack_0, ack => testConfigure_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	249 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_Update/ca
      -- 
    ca_252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_96_inst_ack_1, ack => testConfigure_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	249 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	31 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_final_index_sum_regn_sample_complete
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_final_index_sum_regn_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_final_index_sum_regn_Sample/ack
      -- 
    ack_278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_102_index_offset_ack_0, ack => testConfigure_CP_0_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	249 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (11) 
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_final_index_sum_regn_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_final_index_sum_regn_Update/ack
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_request/$entry
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_request/req
      -- 
    ack_283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_102_index_offset_ack_1, ack => testConfigure_CP_0_elements(18)); -- 
    req_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(18), ack => addr_of_103_final_reg_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_request/$exit
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_request/ack
      -- 
    ack_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_103_final_reg_ack_0, ack => testConfigure_CP_0_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	249 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (28) 
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_complete/ack
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_base_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_word_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_root_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_base_address_resized
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_base_addr_resize/$entry
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_base_addr_resize/$exit
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_base_addr_resize/base_resize_req
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_base_addr_resize/base_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_base_plus_offset/$entry
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_base_plus_offset/$exit
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_base_plus_offset/sum_rename_req
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_base_plus_offset/sum_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_word_addrgen/$entry
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_word_addrgen/$exit
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_word_addrgen/root_register_req
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_word_addrgen/root_register_ack
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/ptr_deref_106_Split/$entry
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/ptr_deref_106_Split/$exit
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/ptr_deref_106_Split/split_req
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/ptr_deref_106_Split/split_ack
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/word_access_start/$entry
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/word_access_start/word_0/$entry
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/word_access_start/word_0/rr
      -- 
    ack_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_103_final_reg_ack_1, ack => testConfigure_CP_0_elements(20)); -- 
    rr_336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(20), ack => ptr_deref_106_store_0_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	30 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Sample/word_access_start/word_0/ra
      -- 
    ra_337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_106_store_0_ack_0, ack => testConfigure_CP_0_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	249 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	31 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Update/word_access_complete/word_0/ca
      -- 
    ca_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_106_store_0_ack_1, ack => testConfigure_CP_0_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	249 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Sample/word_access_start/$entry
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Sample/word_access_start/word_0/rr
      -- 
    rr_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(23), ack => ptr_deref_123_load_0_req_0); -- 
    testConfigure_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(30) & testConfigure_CP_0_elements(249);
      gj_testConfigure_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Sample/word_access_start/$exit
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Sample/word_access_start/word_0/ra
      -- 
    ra_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_123_load_0_ack_0, ack => testConfigure_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	249 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	31 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/word_access_complete/$exit
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/ptr_deref_123_Merge/$entry
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/ptr_deref_123_Merge/$exit
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/ptr_deref_123_Merge/merge_req
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/ptr_deref_123_Merge/merge_ack
      -- 
    ca_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_123_load_0_ack_1, ack => testConfigure_CP_0_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	249 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_update_start_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_Update/cr
      -- 
    ra_407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_131_inst_ack_0, ack => testConfigure_CP_0_elements(26)); -- 
    cr_411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(26), ack => RPIPE_ConvTranspose_input_pipe_131_inst_req_1); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_Sample/rr
      -- 
    ca_412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_131_inst_ack_1, ack => testConfigure_CP_0_elements(27)); -- 
    rr_420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(27), ack => type_cast_135_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_Sample/ra
      -- 
    ra_421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_135_inst_ack_0, ack => testConfigure_CP_0_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	249 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_Update/ca
      -- 
    ca_426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_135_inst_ack_1, ack => testConfigure_CP_0_elements(29)); -- 
    -- CP-element group 30:  transition  delay-element  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	21 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	23 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_ptr_deref_123_delay
      -- 
    -- Element group testConfigure_CP_0_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(21), ack => testConfigure_CP_0_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  branch  join  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	17 
    -- CP-element group 31: 	22 
    -- CP-element group 31: 	25 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (10) 
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136__exit__
      -- CP-element group 31: 	 branch_block_stmt_33/if_stmt_137__entry__
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/$exit
      -- CP-element group 31: 	 branch_block_stmt_33/if_stmt_137_dead_link/$entry
      -- CP-element group 31: 	 branch_block_stmt_33/if_stmt_137_eval_test/$entry
      -- CP-element group 31: 	 branch_block_stmt_33/if_stmt_137_eval_test/$exit
      -- CP-element group 31: 	 branch_block_stmt_33/if_stmt_137_eval_test/branch_req
      -- CP-element group 31: 	 branch_block_stmt_33/R_cmp_138_place
      -- CP-element group 31: 	 branch_block_stmt_33/if_stmt_137_if_link/$entry
      -- CP-element group 31: 	 branch_block_stmt_33/if_stmt_137_else_link/$entry
      -- 
    branch_req_435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(31), ack => if_stmt_137_branch_req_0); -- 
    testConfigure_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(16) & testConfigure_CP_0_elements(17) & testConfigure_CP_0_elements(22) & testConfigure_CP_0_elements(25) & testConfigure_CP_0_elements(29);
      gj_testConfigure_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  place  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	234 
    -- CP-element group 32: 	235 
    -- CP-element group 32: 	237 
    -- CP-element group 32: 	238 
    -- CP-element group 32:  members (20) 
      -- CP-element group 32: 	 branch_block_stmt_33/if_stmt_137_if_link/$exit
      -- CP-element group 32: 	 branch_block_stmt_33/if_stmt_137_if_link/if_choice_transition
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/SplitProtocol/Update/cr
      -- 
    if_choice_transition_440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_137_branch_ack_1, ack => testConfigure_CP_0_elements(32)); -- 
    rr_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_77_inst_req_0); -- 
    cr_2668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_77_inst_req_1); -- 
    rr_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_84_inst_req_0); -- 
    cr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_84_inst_req_1); -- 
    -- CP-element group 33:  fork  transition  place  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	250 
    -- CP-element group 33: 	251 
    -- CP-element group 33:  members (12) 
      -- CP-element group 33: 	 branch_block_stmt_33/if_stmt_137_else_link/$exit
      -- CP-element group 33: 	 branch_block_stmt_33/if_stmt_137_else_link/else_choice_transition
      -- CP-element group 33: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 33: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/SplitProtocol/Update/cr
      -- 
    else_choice_transition_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_137_branch_ack_0, ack => testConfigure_CP_0_elements(33)); -- 
    rr_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => type_cast_147_inst_req_0); -- 
    cr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => type_cast_147_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	261 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/word_access_start/$exit
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/word_access_start/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/word_access_start/word_0/ra
      -- 
    ra_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_165_store_0_ack_0, ack => testConfigure_CP_0_elements(34)); -- 
    -- CP-element group 35:  branch  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	261 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (15) 
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173__exit__
      -- CP-element group 35: 	 branch_block_stmt_33/if_stmt_174__entry__
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/$exit
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Update/word_access_complete/$exit
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Update/word_access_complete/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Update/word_access_complete/word_0/ca
      -- CP-element group 35: 	 branch_block_stmt_33/if_stmt_174_dead_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_33/if_stmt_174_eval_test/$entry
      -- CP-element group 35: 	 branch_block_stmt_33/if_stmt_174_eval_test/$exit
      -- CP-element group 35: 	 branch_block_stmt_33/if_stmt_174_eval_test/branch_req
      -- CP-element group 35: 	 branch_block_stmt_33/R_cmp12223_175_place
      -- CP-element group 35: 	 branch_block_stmt_33/if_stmt_174_if_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_33/if_stmt_174_else_link/$entry
      -- 
    ca_499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_165_store_0_ack_1, ack => testConfigure_CP_0_elements(35)); -- 
    branch_req_507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(35), ack => if_stmt_174_branch_req_0); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	268 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_33/if_stmt_174_if_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_33/if_stmt_174_if_link/if_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_33/forx_xend_bbx_xnph221
      -- CP-element group 36: 	 branch_block_stmt_33/forx_xend_bbx_xnph221_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_33/forx_xend_bbx_xnph221_PhiReq/$exit
      -- 
    if_choice_transition_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_174_branch_ack_1, ack => testConfigure_CP_0_elements(36)); -- 
    -- CP-element group 37:  merge  transition  place  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	265 
    -- CP-element group 37:  members (14) 
      -- CP-element group 37: 	 branch_block_stmt_33/merge_stmt_180__exit__
      -- CP-element group 37: 	 branch_block_stmt_33/forx_xbody14x_xpreheader_forx_xbody14
      -- CP-element group 37: 	 branch_block_stmt_33/if_stmt_174_else_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_33/if_stmt_174_else_link/else_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_33/forx_xend_forx_xbody14x_xpreheader
      -- CP-element group 37: 	 branch_block_stmt_33/forx_xend_forx_xbody14x_xpreheader_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_33/forx_xend_forx_xbody14x_xpreheader_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_33/merge_stmt_180_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_33/merge_stmt_180_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_33/merge_stmt_180_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_33/merge_stmt_180_PhiAck/dummy
      -- CP-element group 37: 	 branch_block_stmt_33/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_33/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_183/$entry
      -- CP-element group 37: 	 branch_block_stmt_33/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/$entry
      -- 
    else_choice_transition_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_174_branch_ack_0, ack => testConfigure_CP_0_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	267 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_Sample/ra
      -- 
    ra_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_199_inst_ack_0, ack => testConfigure_CP_0_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	267 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	55 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_Update/ca
      -- 
    ca_535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_199_inst_ack_1, ack => testConfigure_CP_0_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	267 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	55 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_final_index_sum_regn_sample_complete
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_final_index_sum_regn_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_final_index_sum_regn_Sample/ack
      -- 
    ack_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_205_index_offset_ack_0, ack => testConfigure_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	267 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (11) 
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_offset_calculated
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_final_index_sum_regn_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_final_index_sum_regn_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_request/$entry
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_request/req
      -- 
    ack_566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_205_index_offset_ack_1, ack => testConfigure_CP_0_elements(41)); -- 
    req_575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(41), ack => addr_of_206_final_reg_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_request/$exit
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_request/ack
      -- 
    ack_576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_206_final_reg_ack_0, ack => testConfigure_CP_0_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	267 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	48 
    -- CP-element group 43:  members (19) 
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_complete/ack
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_base_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_word_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_root_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_base_address_resized
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_base_addr_resize/$entry
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_base_addr_resize/$exit
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_base_addr_resize/base_resize_req
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_base_addr_resize/base_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_base_plus_offset/$entry
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_base_plus_offset/$exit
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_base_plus_offset/sum_rename_req
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_base_plus_offset/sum_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_word_addrgen/$entry
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_word_addrgen/$exit
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_word_addrgen/root_register_req
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_word_addrgen/root_register_ack
      -- 
    ack_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_206_final_reg_ack_1, ack => testConfigure_CP_0_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	267 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_update_start_
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_Update/cr
      -- 
    ra_590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_209_inst_ack_0, ack => testConfigure_CP_0_elements(44)); -- 
    cr_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(44), ack => RPIPE_ConvTranspose_input_pipe_209_inst_req_1); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_Sample/rr
      -- 
    ca_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_209_inst_ack_1, ack => testConfigure_CP_0_elements(45)); -- 
    rr_603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(45), ack => type_cast_213_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_Sample/ra
      -- 
    ra_604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_213_inst_ack_0, ack => testConfigure_CP_0_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	267 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_Update/ca
      -- 
    ca_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_213_inst_ack_1, ack => testConfigure_CP_0_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	43 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/ptr_deref_216_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/ptr_deref_216_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/ptr_deref_216_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/ptr_deref_216_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/word_access_start/word_0/rr
      -- 
    rr_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(48), ack => ptr_deref_216_store_0_req_0); -- 
    testConfigure_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(47) & testConfigure_CP_0_elements(43);
      gj_testConfigure_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	54 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Sample/word_access_start/word_0/ra
      -- 
    ra_648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_216_store_0_ack_0, ack => testConfigure_CP_0_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	267 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	55 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Update/word_access_complete/word_0/ca
      -- 
    ca_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_216_store_0_ack_1, ack => testConfigure_CP_0_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: 	267 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Sample/word_access_start/word_0/rr
      -- 
    rr_692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(51), ack => ptr_deref_233_load_0_req_0); -- 
    testConfigure_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(54) & testConfigure_CP_0_elements(267);
      gj_testConfigure_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Sample/word_access_start/word_0/ra
      -- 
    ra_693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_233_load_0_ack_0, ack => testConfigure_CP_0_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	267 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/word_access_complete/word_0/ca
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/ptr_deref_233_Merge/$entry
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/ptr_deref_233_Merge/$exit
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/ptr_deref_233_Merge/merge_req
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/ptr_deref_233_Merge/merge_ack
      -- 
    ca_704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_233_load_0_ack_1, ack => testConfigure_CP_0_elements(53)); -- 
    -- CP-element group 54:  transition  delay-element  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	49 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_ptr_deref_233_delay
      -- 
    -- Element group testConfigure_CP_0_elements(54) is a control-delay.
    cp_element_54_delay: control_delay_element  generic map(name => " 54_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(49), ack => testConfigure_CP_0_elements(54), clk => clk, reset =>reset);
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	50 
    -- CP-element group 55: 	39 
    -- CP-element group 55: 	40 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239__exit__
      -- CP-element group 55: 	 branch_block_stmt_33/if_stmt_240__entry__
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/$exit
      -- CP-element group 55: 	 branch_block_stmt_33/if_stmt_240_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_33/if_stmt_240_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_33/if_stmt_240_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_33/if_stmt_240_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_33/R_cmp12_241_place
      -- CP-element group 55: 	 branch_block_stmt_33/if_stmt_240_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_33/if_stmt_240_else_link/$entry
      -- 
    branch_req_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => if_stmt_240_branch_req_0); -- 
    testConfigure_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(50) & testConfigure_CP_0_elements(39) & testConfigure_CP_0_elements(40) & testConfigure_CP_0_elements(53);
      gj_testConfigure_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	262 
    -- CP-element group 56: 	263 
    -- CP-element group 56:  members (12) 
      -- CP-element group 56: 	 branch_block_stmt_33/if_stmt_240_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_33/if_stmt_240_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14
      -- CP-element group 56: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/$entry
      -- CP-element group 56: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/$entry
      -- CP-element group 56: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/SplitProtocol/Update/cr
      -- 
    if_choice_transition_723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_240_branch_ack_1, ack => testConfigure_CP_0_elements(56)); -- 
    rr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_186_inst_req_0); -- 
    cr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_186_inst_req_1); -- 
    -- CP-element group 57:  merge  transition  place  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	268 
    -- CP-element group 57:  members (13) 
      -- CP-element group 57: 	 branch_block_stmt_33/merge_stmt_246__exit__
      -- CP-element group 57: 	 branch_block_stmt_33/bbx_xnph221x_xloopexit_bbx_xnph221
      -- CP-element group 57: 	 branch_block_stmt_33/if_stmt_240_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_33/if_stmt_240_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_33/forx_xbody14_bbx_xnph221x_xloopexit
      -- CP-element group 57: 	 branch_block_stmt_33/forx_xbody14_bbx_xnph221x_xloopexit_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_33/forx_xbody14_bbx_xnph221x_xloopexit_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_33/merge_stmt_246_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_33/merge_stmt_246_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_33/merge_stmt_246_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_33/merge_stmt_246_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_33/bbx_xnph221x_xloopexit_bbx_xnph221_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_33/bbx_xnph221x_xloopexit_bbx_xnph221_PhiReq/$exit
      -- 
    else_choice_transition_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_240_branch_ack_0, ack => testConfigure_CP_0_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	268 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_update_start_
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_Update/cr
      -- 
    ra_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_250_inst_ack_0, ack => testConfigure_CP_0_elements(58)); -- 
    cr_745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(58), ack => RPIPE_ConvTranspose_input_pipe_250_inst_req_1); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_Sample/rr
      -- 
    ca_746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_250_inst_ack_1, ack => testConfigure_CP_0_elements(59)); -- 
    rr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(59), ack => type_cast_254_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_Sample/ra
      -- 
    ra_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_254_inst_ack_0, ack => testConfigure_CP_0_elements(60)); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	268 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	269 
    -- CP-element group 61: 	270 
    -- CP-element group 61: 	271 
    -- CP-element group 61:  members (17) 
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255__exit__
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/$exit
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_258/$entry
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/$entry
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/$entry
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/SplitProtocol/Update/cr
      -- 
    ca_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_254_inst_ack_1, ack => testConfigure_CP_0_elements(61)); -- 
    rr_2929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(61), ack => type_cast_268_inst_req_0); -- 
    cr_2934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(61), ack => type_cast_268_inst_req_1); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	284 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_request/$exit
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_request/ack
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_sample_completed_
      -- 
    ack_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_275_final_reg_ack_0, ack => testConfigure_CP_0_elements(62)); -- 
    -- CP-element group 63:  join  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	284 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (28) 
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_complete/ack
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_base_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_word_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_root_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_base_address_resized
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_base_addr_resize/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_base_addr_resize/$exit
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_base_addr_resize/base_resize_req
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_base_addr_resize/base_resize_ack
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_base_plus_offset/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_base_plus_offset/$exit
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_base_plus_offset/sum_rename_req
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_base_plus_offset/sum_rename_ack
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_word_addrgen/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_word_addrgen/$exit
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_word_addrgen/root_register_req
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_word_addrgen/root_register_ack
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/ptr_deref_278_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/ptr_deref_278_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/ptr_deref_278_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/ptr_deref_278_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/word_access_start/word_0/rr
      -- 
    ack_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_275_final_reg_ack_1, ack => testConfigure_CP_0_elements(63)); -- 
    rr_840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(63), ack => ptr_deref_278_store_0_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Sample/word_access_start/word_0/ra
      -- 
    ra_841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_278_store_0_ack_0, ack => testConfigure_CP_0_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	284 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	70 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Update/word_access_complete/word_0/ca
      -- 
    ca_852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_278_store_0_ack_1, ack => testConfigure_CP_0_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	284 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_update_start_
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_Update/cr
      -- 
    ra_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_282_inst_ack_0, ack => testConfigure_CP_0_elements(66)); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(66), ack => RPIPE_ConvTranspose_input_pipe_282_inst_req_1); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_Sample/rr
      -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_282_inst_ack_1, ack => testConfigure_CP_0_elements(67)); -- 
    rr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(67), ack => type_cast_286_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_Sample/ra
      -- 
    ra_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_286_inst_ack_0, ack => testConfigure_CP_0_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	284 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_Update/ca
      -- 
    ca_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_286_inst_ack_1, ack => testConfigure_CP_0_elements(69)); -- 
    -- CP-element group 70:  branch  join  transition  place  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	65 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (10) 
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299__exit__
      -- CP-element group 70: 	 branch_block_stmt_33/if_stmt_300__entry__
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/$exit
      -- CP-element group 70: 	 branch_block_stmt_33/if_stmt_300_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_33/if_stmt_300_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_33/if_stmt_300_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_33/if_stmt_300_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_33/R_exitcond_301_place
      -- CP-element group 70: 	 branch_block_stmt_33/if_stmt_300_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_33/if_stmt_300_else_link/$entry
      -- 
    branch_req_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(70), ack => if_stmt_300_branch_req_0); -- 
    testConfigure_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(65) & testConfigure_CP_0_elements(69);
      gj_testConfigure_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	285 
    -- CP-element group 71: 	286 
    -- CP-element group 71:  members (12) 
      -- CP-element group 71: 	 branch_block_stmt_33/if_stmt_300_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_33/if_stmt_300_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_33/forx_xbody28_forx_xend37
      -- CP-element group 71: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/$entry
      -- CP-element group 71: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/$entry
      -- CP-element group 71: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/$entry
      -- CP-element group 71: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/SplitProtocol/$entry
      -- CP-element group 71: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/SplitProtocol/Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/SplitProtocol/Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/SplitProtocol/Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/SplitProtocol/Update/cr
      -- 
    if_choice_transition_893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_300_branch_ack_1, ack => testConfigure_CP_0_elements(71)); -- 
    rr_3014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(71), ack => type_cast_310_inst_req_0); -- 
    cr_3019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(71), ack => type_cast_310_inst_req_1); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	274 
    -- CP-element group 72: 	275 
    -- CP-element group 72: 	277 
    -- CP-element group 72: 	278 
    -- CP-element group 72:  members (20) 
      -- CP-element group 72: 	 branch_block_stmt_33/if_stmt_300_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_33/if_stmt_300_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/SplitProtocol/Update/cr
      -- 
    else_choice_transition_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_300_branch_ack_0, ack => testConfigure_CP_0_elements(72)); -- 
    rr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_264_inst_req_0); -- 
    cr_2960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_264_inst_req_1); -- 
    rr_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_270_inst_req_0); -- 
    cr_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_270_inst_req_1); -- 
    -- CP-element group 73:  join  fork  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	288 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: 	75 
    -- CP-element group 73: 	76 
    -- CP-element group 73: 	79 
    -- CP-element group 73: 	80 
    -- CP-element group 73: 	82 
    -- CP-element group 73: 	86 
    -- CP-element group 73: 	87 
    -- CP-element group 73: 	89 
    -- CP-element group 73: 	93 
    -- CP-element group 73: 	94 
    -- CP-element group 73: 	96 
    -- CP-element group 73: 	97 
    -- CP-element group 73: 	98 
    -- CP-element group 73: 	99 
    -- CP-element group 73: 	100 
    -- CP-element group 73: 	101 
    -- CP-element group 73: 	102 
    -- CP-element group 73: 	105 
    -- CP-element group 73: 	106 
    -- CP-element group 73: 	107 
    -- CP-element group 73: 	108 
    -- CP-element group 73: 	109 
    -- CP-element group 73: 	110 
    -- CP-element group 73: 	111 
    -- CP-element group 73: 	112 
    -- CP-element group 73: 	113 
    -- CP-element group 73: 	116 
    -- CP-element group 73:  members (280) 
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/STORE_padding_312_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/STORE_padding_312_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/STORE_padding_312_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/STORE_padding_312_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_update_start_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Update/word_access_complete/word_0/cr
      -- 
    cr_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => STORE_padding_312_store_0_req_1); -- 
    rr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => STORE_padding_312_store_0_req_0); -- 
    rr_943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_0); -- 
    cr_962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_320_inst_req_1); -- 
    cr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_331_store_0_req_1); -- 
    cr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_339_inst_req_1); -- 
    cr_1090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_350_store_0_req_1); -- 
    cr_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_358_inst_req_1); -- 
    cr_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_369_store_0_req_1); -- 
    cr_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_382_load_0_req_1); -- 
    rr_1202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_382_load_0_req_0); -- 
    cr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_394_load_0_req_1); -- 
    rr_1252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_394_load_0_req_0); -- 
    cr_1313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_406_load_0_req_1); -- 
    rr_1302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_406_load_0_req_0); -- 
    cr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_420_inst_req_1); -- 
    cr_1377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_432_load_0_req_1); -- 
    rr_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_432_load_0_req_0); -- 
    cr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_444_load_0_req_1); -- 
    rr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_444_load_0_req_0); -- 
    cr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_456_load_0_req_1); -- 
    rr_1466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_456_load_0_req_0); -- 
    cr_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_468_load_0_req_1); -- 
    rr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_468_load_0_req_0); -- 
    cr_1546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_487_inst_req_1); -- 
    testConfigure_CP_0_elements(73) <= testConfigure_CP_0_elements(288);
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Sample/word_access_start/word_0/ra
      -- 
    ra_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_312_store_0_ack_0, ack => testConfigure_CP_0_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	119 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/STORE_padding_312_Update/word_access_complete/word_0/ca
      -- 
    ca_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_312_store_0_ack_1, ack => testConfigure_CP_0_elements(75)); -- 
    -- CP-element group 76:  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	73 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_update_start_
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_Update/cr
      -- 
    ra_944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_0, ack => testConfigure_CP_0_elements(76)); -- 
    cr_948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_1); -- 
    -- CP-element group 77:  fork  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	83 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_316_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_Sample/rr
      -- 
    ca_949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_1, ack => testConfigure_CP_0_elements(77)); -- 
    rr_957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_320_inst_req_0); -- 
    rr_1021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => RPIPE_ConvTranspose_input_pipe_335_inst_req_0); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_Sample/ra
      -- 
    ra_958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_0, ack => testConfigure_CP_0_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	73 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_320_Update/ca
      -- 
    ca_963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_1, ack => testConfigure_CP_0_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	73 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/ptr_deref_331_Split/$entry
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/ptr_deref_331_Split/$exit
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/ptr_deref_331_Split/split_req
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/ptr_deref_331_Split/split_ack
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/word_access_start/$entry
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/word_access_start/word_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/word_access_start/word_0/rr
      -- 
    rr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(80), ack => ptr_deref_331_store_0_req_0); -- 
    testConfigure_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(79);
      gj_testConfigure_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	117 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/word_access_start/$exit
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/word_access_start/word_0/$exit
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Sample/word_access_start/word_0/ra
      -- 
    ra_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_331_store_0_ack_0, ack => testConfigure_CP_0_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	73 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	119 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Update/word_access_complete/$exit
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Update/word_access_complete/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_Update/word_access_complete/word_0/ca
      -- 
    ca_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_331_store_0_ack_1, ack => testConfigure_CP_0_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	77 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_update_start_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_Sample/ra
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_Update/cr
      -- 
    ra_1022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_335_inst_ack_0, ack => testConfigure_CP_0_elements(83)); -- 
    cr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(83), ack => RPIPE_ConvTranspose_input_pipe_335_inst_req_1); -- 
    -- CP-element group 84:  fork  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	90 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_335_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_Sample/rr
      -- 
    ca_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_335_inst_ack_1, ack => testConfigure_CP_0_elements(84)); -- 
    rr_1035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => type_cast_339_inst_req_0); -- 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => RPIPE_ConvTranspose_input_pipe_354_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_Sample/ra
      -- 
    ra_1036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_339_inst_ack_0, ack => testConfigure_CP_0_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	73 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_339_Update/ca
      -- 
    ca_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_339_inst_ack_1, ack => testConfigure_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	73 
    -- CP-element group 87: 	86 
    -- CP-element group 87: 	117 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/ptr_deref_350_Split/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/ptr_deref_350_Split/$exit
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/ptr_deref_350_Split/split_req
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/ptr_deref_350_Split/split_ack
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/word_access_start/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/word_access_start/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/word_access_start/word_0/rr
      -- 
    rr_1079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(87), ack => ptr_deref_350_store_0_req_0); -- 
    testConfigure_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(86) & testConfigure_CP_0_elements(117);
      gj_testConfigure_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	118 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/word_access_start/$exit
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/word_access_start/word_0/$exit
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Sample/word_access_start/word_0/ra
      -- 
    ra_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_350_store_0_ack_0, ack => testConfigure_CP_0_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	73 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	119 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Update/word_access_complete/$exit
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Update/word_access_complete/word_0/$exit
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_Update/word_access_complete/word_0/ca
      -- 
    ca_1091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_350_store_0_ack_1, ack => testConfigure_CP_0_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	84 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_update_start_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_Update/cr
      -- 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_354_inst_ack_0, ack => testConfigure_CP_0_elements(90)); -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(90), ack => RPIPE_ConvTranspose_input_pipe_354_inst_req_1); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/RPIPE_ConvTranspose_input_pipe_354_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_sample_start_
      -- 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_354_inst_ack_1, ack => testConfigure_CP_0_elements(91)); -- 
    rr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(91), ack => type_cast_358_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_sample_completed_
      -- 
    ra_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_0, ack => testConfigure_CP_0_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	73 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_Update/ca
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_358_Update/$exit
      -- 
    ca_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_1, ack => testConfigure_CP_0_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	73 
    -- CP-element group 94: 	93 
    -- CP-element group 94: 	118 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/word_access_start/word_0/rr
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/word_access_start/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/word_access_start/$entry
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/ptr_deref_369_Split/split_ack
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/ptr_deref_369_Split/split_req
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/ptr_deref_369_Split/$exit
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/ptr_deref_369_Split/$entry
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/$entry
      -- 
    rr_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(94), ack => ptr_deref_369_store_0_req_0); -- 
    testConfigure_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(93) & testConfigure_CP_0_elements(118);
      gj_testConfigure_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/word_access_start/word_0/ra
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/word_access_start/word_0/$exit
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/word_access_start/$exit
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Sample/$exit
      -- 
    ra_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_369_store_0_ack_0, ack => testConfigure_CP_0_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	73 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	119 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Update/word_access_complete/$exit
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Update/word_access_complete/word_0/ca
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_369_Update/word_access_complete/word_0/$exit
      -- 
    ca_1169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_369_store_0_ack_1, ack => testConfigure_CP_0_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	73 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Sample/word_access_start/word_0/ra
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Sample/word_access_start/word_0/$exit
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Sample/word_access_start/$exit
      -- 
    ra_1203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_382_load_0_ack_0, ack => testConfigure_CP_0_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	73 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	103 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/ptr_deref_382_Merge/merge_ack
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/ptr_deref_382_Merge/merge_req
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/ptr_deref_382_Merge/$exit
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/ptr_deref_382_Merge/$entry
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/word_access_complete/word_0/ca
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/word_access_complete/word_0/$exit
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/word_access_complete/$exit
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_382_update_completed_
      -- 
    ca_1214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_382_load_0_ack_1, ack => testConfigure_CP_0_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	73 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Sample/word_access_start/word_0/ra
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Sample/word_access_start/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Sample/word_access_start/$exit
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Sample/$exit
      -- 
    ra_1253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_394_load_0_ack_0, ack => testConfigure_CP_0_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	73 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/word_access_complete/word_0/$exit
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/word_access_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/ptr_deref_394_Merge/merge_ack
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/ptr_deref_394_Merge/merge_req
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/ptr_deref_394_Merge/$exit
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/ptr_deref_394_Merge/$entry
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_394_Update/word_access_complete/word_0/ca
      -- 
    ca_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_394_load_0_ack_1, ack => testConfigure_CP_0_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	73 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Sample/word_access_start/word_0/ra
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Sample/word_access_start/word_0/$exit
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Sample/word_access_start/$exit
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Sample/$exit
      -- 
    ra_1303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_406_load_0_ack_0, ack => testConfigure_CP_0_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	73 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (9) 
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/ptr_deref_406_Merge/$exit
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/ptr_deref_406_Merge/$entry
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/word_access_complete/word_0/ca
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/word_access_complete/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/word_access_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/ptr_deref_406_Merge/merge_ack
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_406_Update/ptr_deref_406_Merge/merge_req
      -- 
    ca_1314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_406_load_0_ack_1, ack => testConfigure_CP_0_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	98 
    -- CP-element group 103: 	100 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_sample_start_
      -- 
    rr_1327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(103), ack => type_cast_420_inst_req_0); -- 
    testConfigure_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(98) & testConfigure_CP_0_elements(100) & testConfigure_CP_0_elements(102);
      gj_testConfigure_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_sample_completed_
      -- 
    ra_1328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_420_inst_ack_0, ack => testConfigure_CP_0_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	73 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	119 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_420_update_completed_
      -- 
    ca_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_420_inst_ack_1, ack => testConfigure_CP_0_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	73 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Sample/word_access_start/word_0/$exit
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Sample/word_access_start/$exit
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Sample/word_access_start/word_0/ra
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Sample/$exit
      -- 
    ra_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_432_load_0_ack_0, ack => testConfigure_CP_0_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	73 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	114 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/ptr_deref_432_Merge/merge_ack
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/ptr_deref_432_Merge/merge_req
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/ptr_deref_432_Merge/$exit
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/ptr_deref_432_Merge/$entry
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/word_access_complete/word_0/ca
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/word_access_complete/word_0/$exit
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/word_access_complete/$exit
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_432_Update/$exit
      -- 
    ca_1378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_432_load_0_ack_1, ack => testConfigure_CP_0_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	73 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Sample/word_access_start/word_0/ra
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Sample/word_access_start/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Sample/word_access_start/$exit
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Sample/$exit
      -- 
    ra_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_444_load_0_ack_0, ack => testConfigure_CP_0_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	73 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	114 
    -- CP-element group 109:  members (9) 
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/ptr_deref_444_Merge/$exit
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/ptr_deref_444_Merge/merge_req
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/ptr_deref_444_Merge/$entry
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/word_access_complete/word_0/ca
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/word_access_complete/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/word_access_complete/$exit
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_444_Update/ptr_deref_444_Merge/merge_ack
      -- 
    ca_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_444_load_0_ack_1, ack => testConfigure_CP_0_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	73 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Sample/word_access_start/word_0/ra
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Sample/word_access_start/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Sample/word_access_start/$exit
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Sample/$exit
      -- 
    ra_1467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_456_load_0_ack_0, ack => testConfigure_CP_0_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	73 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/word_access_complete/word_0/ca
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/word_access_complete/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/word_access_complete/$exit
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/ptr_deref_456_Merge/merge_ack
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/ptr_deref_456_Merge/merge_req
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/ptr_deref_456_Merge/$exit
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_456_Update/ptr_deref_456_Merge/$entry
      -- 
    ca_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_456_load_0_ack_1, ack => testConfigure_CP_0_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	73 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Sample/word_access_start/word_0/ra
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Sample/word_access_start/word_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Sample/word_access_start/$exit
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Sample/$exit
      -- 
    ra_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_468_load_0_ack_0, ack => testConfigure_CP_0_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	73 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (9) 
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/word_access_complete/$exit
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/word_access_complete/word_0/ca
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/ptr_deref_468_Merge/merge_req
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/ptr_deref_468_Merge/$entry
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/ptr_deref_468_Merge/$exit
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/word_access_complete/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_Update/ptr_deref_468_Merge/merge_ack
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_468_update_completed_
      -- 
    ca_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_468_load_0_ack_1, ack => testConfigure_CP_0_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	107 
    -- CP-element group 114: 	109 
    -- CP-element group 114: 	111 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_sample_start_
      -- 
    rr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(114), ack => type_cast_487_inst_req_0); -- 
    testConfigure_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(107) & testConfigure_CP_0_elements(109) & testConfigure_CP_0_elements(111) & testConfigure_CP_0_elements(113);
      gj_testConfigure_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_sample_completed_
      -- 
    ra_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_487_inst_ack_0, ack => testConfigure_CP_0_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	73 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/type_cast_487_update_completed_
      -- 
    ca_1547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_487_inst_ack_1, ack => testConfigure_CP_0_elements(116)); -- 
    -- CP-element group 117:  transition  delay-element  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	81 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	87 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_331_ptr_deref_350_delay
      -- 
    -- Element group testConfigure_CP_0_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(81), ack => testConfigure_CP_0_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  transition  delay-element  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	88 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	94 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/ptr_deref_350_ptr_deref_369_delay
      -- 
    -- Element group testConfigure_CP_0_elements(118) is a control-delay.
    cp_element_118_delay: control_delay_element  generic map(name => " 118_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(88), ack => testConfigure_CP_0_elements(118), clk => clk, reset =>reset);
    -- CP-element group 119:  branch  join  transition  place  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	75 
    -- CP-element group 119: 	82 
    -- CP-element group 119: 	89 
    -- CP-element group 119: 	96 
    -- CP-element group 119: 	105 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (10) 
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_501_else_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_501_eval_test/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_501_eval_test/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_501_dead_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_501_eval_test/branch_req
      -- CP-element group 119: 	 branch_block_stmt_33/R_cmp65213_502_place
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_501_if_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500__exit__
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_501__entry__
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500/$exit
      -- 
    branch_req_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => if_stmt_501_branch_req_0); -- 
    testConfigure_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(75) & testConfigure_CP_0_elements(82) & testConfigure_CP_0_elements(89) & testConfigure_CP_0_elements(96) & testConfigure_CP_0_elements(105) & testConfigure_CP_0_elements(116);
      gj_testConfigure_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	289 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_33/if_stmt_501_if_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_33/if_stmt_501_if_link/if_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_33/forx_xend37_forx_xcond119x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_33/forx_xend37_forx_xcond119x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_33/forx_xend37_forx_xcond119x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_501_branch_ack_1, ack => testConfigure_CP_0_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	124 
    -- CP-element group 121: 	125 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_33/if_stmt_501_else_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/if_stmt_501_else_link/else_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_528__exit__
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561__entry__
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xend37_bbx_xnph215
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_update_start_
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xend37_bbx_xnph215_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xend37_bbx_xnph215_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_528_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_528_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_528_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_528_PhiAck/dummy
      -- 
    else_choice_transition_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_501_branch_ack_0, ack => testConfigure_CP_0_elements(121)); -- 
    rr_1601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(121), ack => type_cast_541_inst_req_0); -- 
    cr_1606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(121), ack => type_cast_541_inst_req_1); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	289 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	302 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_33/if_stmt_522_if_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_33/if_stmt_522_if_link/if_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond119x_xpreheader_forx_xend180
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond119x_xpreheader_forx_xend180_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond119x_xpreheader_forx_xend180_PhiReq/$exit
      -- 
    if_choice_transition_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_522_branch_ack_1, ack => testConfigure_CP_0_elements(122)); -- 
    -- CP-element group 123:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	289 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	168 
    -- CP-element group 123: 	169 
    -- CP-element group 123:  members (18) 
      -- CP-element group 123: 	 branch_block_stmt_33/merge_stmt_733__exit__
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771__entry__
      -- CP-element group 123: 	 branch_block_stmt_33/if_stmt_522_else_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_33/if_stmt_522_else_link/else_choice_transition
      -- CP-element group 123: 	 branch_block_stmt_33/forx_xcond119x_xpreheader_bbx_xnph210
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/$entry
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_update_start_
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_Update/cr
      -- CP-element group 123: 	 branch_block_stmt_33/forx_xcond119x_xpreheader_bbx_xnph210_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_33/forx_xcond119x_xpreheader_bbx_xnph210_PhiReq/$exit
      -- CP-element group 123: 	 branch_block_stmt_33/merge_stmt_733_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_33/merge_stmt_733_PhiAck/$entry
      -- CP-element group 123: 	 branch_block_stmt_33/merge_stmt_733_PhiAck/$exit
      -- CP-element group 123: 	 branch_block_stmt_33/merge_stmt_733_PhiAck/dummy
      -- 
    else_choice_transition_1588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_522_branch_ack_0, ack => testConfigure_CP_0_elements(123)); -- 
    rr_1960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(123), ack => type_cast_751_inst_req_0); -- 
    cr_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(123), ack => type_cast_751_inst_req_1); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_Sample/ra
      -- 
    ra_1602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_0, ack => testConfigure_CP_0_elements(124)); -- 
    -- CP-element group 125:  transition  place  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	121 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	290 
    -- CP-element group 125:  members (9) 
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561__exit__
      -- CP-element group 125: 	 branch_block_stmt_33/bbx_xnph215_forx_xbody67
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/$exit
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_533_to_assign_stmt_561/type_cast_541_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_33/bbx_xnph215_forx_xbody67_PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_33/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_564/$entry
      -- CP-element group 125: 	 branch_block_stmt_33/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/$entry
      -- 
    ca_1607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_1, ack => testConfigure_CP_0_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	295 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	165 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_final_index_sum_regn_sample_complete
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_final_index_sum_regn_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_final_index_sum_regn_Sample/ack
      -- 
    ack_1636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_576_index_offset_ack_0, ack => testConfigure_CP_0_elements(126)); -- 
    -- CP-element group 127:  transition  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	295 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (11) 
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_root_address_calculated
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_offset_calculated
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_final_index_sum_regn_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_final_index_sum_regn_Update/ack
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_base_plus_offset/$entry
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_base_plus_offset/$exit
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_base_plus_offset/sum_rename_req
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_base_plus_offset/sum_rename_ack
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_request/$entry
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_request/req
      -- 
    ack_1641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_576_index_offset_ack_1, ack => testConfigure_CP_0_elements(127)); -- 
    req_1650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(127), ack => addr_of_577_final_reg_req_0); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_request/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_request/ack
      -- 
    ack_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_577_final_reg_ack_0, ack => testConfigure_CP_0_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	295 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	162 
    -- CP-element group 129:  members (19) 
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_complete/$exit
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_complete/ack
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_base_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_word_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_root_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_base_address_resized
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_base_addr_resize/$entry
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_base_addr_resize/$exit
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_base_addr_resize/base_resize_req
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_base_addr_resize/base_resize_ack
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_base_plus_offset/$entry
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_base_plus_offset/$exit
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_base_plus_offset/sum_rename_req
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_base_plus_offset/sum_rename_ack
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_word_addrgen/$entry
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_word_addrgen/$exit
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_word_addrgen/root_register_req
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_word_addrgen/root_register_ack
      -- 
    ack_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_577_final_reg_ack_1, ack => testConfigure_CP_0_elements(129)); -- 
    -- CP-element group 130:  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	295 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (6) 
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_update_start_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_Sample/ra
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_Update/cr
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_580_inst_ack_0, ack => testConfigure_CP_0_elements(130)); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(130), ack => RPIPE_ConvTranspose_input_pipe_580_inst_req_1); -- 
    -- CP-element group 131:  fork  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	134 
    -- CP-element group 131:  members (9) 
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_Sample/rr
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_580_inst_ack_1, ack => testConfigure_CP_0_elements(131)); -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => type_cast_584_inst_req_0); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => RPIPE_ConvTranspose_input_pipe_593_inst_req_0); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_Sample/ra
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_584_inst_ack_0, ack => testConfigure_CP_0_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	295 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	162 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_Update/ca
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_584_inst_ack_1, ack => testConfigure_CP_0_elements(133)); -- 
    -- CP-element group 134:  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	131 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_update_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_Sample/ra
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_Update/cr
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_593_inst_ack_0, ack => testConfigure_CP_0_elements(134)); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(134), ack => RPIPE_ConvTranspose_input_pipe_593_inst_req_1); -- 
    -- CP-element group 135:  fork  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: 	138 
    -- CP-element group 135:  members (9) 
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_593_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_Sample/rr
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_Sample/rr
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_593_inst_ack_1, ack => testConfigure_CP_0_elements(135)); -- 
    rr_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(135), ack => type_cast_597_inst_req_0); -- 
    rr_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(135), ack => RPIPE_ConvTranspose_input_pipe_611_inst_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_Sample/ra
      -- 
    ra_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_597_inst_ack_0, ack => testConfigure_CP_0_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	295 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	162 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_Update/ca
      -- 
    ca_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_597_inst_ack_1, ack => testConfigure_CP_0_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_update_start_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_Update/cr
      -- 
    ra_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_611_inst_ack_0, ack => testConfigure_CP_0_elements(138)); -- 
    cr_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(138), ack => RPIPE_ConvTranspose_input_pipe_611_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	142 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_611_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_Sample/rr
      -- 
    ca_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_611_inst_ack_1, ack => testConfigure_CP_0_elements(139)); -- 
    rr_1734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => type_cast_615_inst_req_0); -- 
    rr_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => RPIPE_ConvTranspose_input_pipe_629_inst_req_0); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_Sample/ra
      -- 
    ra_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_0, ack => testConfigure_CP_0_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	295 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	162 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_Update/ca
      -- 
    ca_1740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_1, ack => testConfigure_CP_0_elements(141)); -- 
    -- CP-element group 142:  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (6) 
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_update_start_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_Sample/ra
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_Update/cr
      -- 
    ra_1749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_629_inst_ack_0, ack => testConfigure_CP_0_elements(142)); -- 
    cr_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(142), ack => RPIPE_ConvTranspose_input_pipe_629_inst_req_1); -- 
    -- CP-element group 143:  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143: 	146 
    -- CP-element group 143:  members (9) 
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_629_Update/ca
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_Sample/rr
      -- 
    ca_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_629_inst_ack_1, ack => testConfigure_CP_0_elements(143)); -- 
    rr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => type_cast_633_inst_req_0); -- 
    rr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => RPIPE_ConvTranspose_input_pipe_647_inst_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_Sample/ra
      -- 
    ra_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_633_inst_ack_0, ack => testConfigure_CP_0_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	295 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	162 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_Update/ca
      -- 
    ca_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_633_inst_ack_1, ack => testConfigure_CP_0_elements(145)); -- 
    -- CP-element group 146:  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	143 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (6) 
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_update_start_
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_Update/cr
      -- 
    ra_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_647_inst_ack_0, ack => testConfigure_CP_0_elements(146)); -- 
    cr_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(146), ack => RPIPE_ConvTranspose_input_pipe_647_inst_req_1); -- 
    -- CP-element group 147:  fork  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147: 	150 
    -- CP-element group 147:  members (9) 
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_647_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_Sample/rr
      -- 
    ca_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_647_inst_ack_1, ack => testConfigure_CP_0_elements(147)); -- 
    rr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => type_cast_651_inst_req_0); -- 
    rr_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => RPIPE_ConvTranspose_input_pipe_665_inst_req_0); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_Sample/ra
      -- 
    ra_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_651_inst_ack_0, ack => testConfigure_CP_0_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	295 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	162 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_Update/ca
      -- 
    ca_1796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_651_inst_ack_1, ack => testConfigure_CP_0_elements(149)); -- 
    -- CP-element group 150:  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	147 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (6) 
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_update_start_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_Update/cr
      -- 
    ra_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_665_inst_ack_0, ack => testConfigure_CP_0_elements(150)); -- 
    cr_1809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(150), ack => RPIPE_ConvTranspose_input_pipe_665_inst_req_1); -- 
    -- CP-element group 151:  fork  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: 	154 
    -- CP-element group 151:  members (9) 
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_665_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_Sample/rr
      -- 
    ca_1810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_665_inst_ack_1, ack => testConfigure_CP_0_elements(151)); -- 
    rr_1818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => type_cast_669_inst_req_0); -- 
    rr_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => RPIPE_ConvTranspose_input_pipe_683_inst_req_0); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_Sample/ra
      -- 
    ra_1819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_669_inst_ack_0, ack => testConfigure_CP_0_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	295 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	162 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_Update/ca
      -- 
    ca_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_669_inst_ack_1, ack => testConfigure_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	151 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_update_start_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_Update/cr
      -- 
    ra_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_683_inst_ack_0, ack => testConfigure_CP_0_elements(154)); -- 
    cr_1837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(154), ack => RPIPE_ConvTranspose_input_pipe_683_inst_req_1); -- 
    -- CP-element group 155:  fork  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	158 
    -- CP-element group 155:  members (9) 
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_683_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_Sample/rr
      -- 
    ca_1838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_683_inst_ack_1, ack => testConfigure_CP_0_elements(155)); -- 
    rr_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => type_cast_687_inst_req_0); -- 
    rr_1860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => RPIPE_ConvTranspose_input_pipe_701_inst_req_0); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_Sample/ra
      -- 
    ra_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_0, ack => testConfigure_CP_0_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	295 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	162 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_Update/ca
      -- 
    ca_1852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_1, ack => testConfigure_CP_0_elements(157)); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	155 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_update_start_
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_Update/cr
      -- 
    ra_1861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_701_inst_ack_0, ack => testConfigure_CP_0_elements(158)); -- 
    cr_1865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(158), ack => RPIPE_ConvTranspose_input_pipe_701_inst_req_1); -- 
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (6) 
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_701_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_Sample/rr
      -- 
    ca_1866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_701_inst_ack_1, ack => testConfigure_CP_0_elements(159)); -- 
    rr_1874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(159), ack => type_cast_705_inst_req_0); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_Sample/ra
      -- 
    ra_1875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_705_inst_ack_0, ack => testConfigure_CP_0_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	295 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_Update/ca
      -- 
    ca_1880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_705_inst_ack_1, ack => testConfigure_CP_0_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	129 
    -- CP-element group 162: 	133 
    -- CP-element group 162: 	137 
    -- CP-element group 162: 	141 
    -- CP-element group 162: 	145 
    -- CP-element group 162: 	149 
    -- CP-element group 162: 	153 
    -- CP-element group 162: 	157 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (9) 
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/ptr_deref_713_Split/$entry
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/ptr_deref_713_Split/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/ptr_deref_713_Split/split_req
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/ptr_deref_713_Split/split_ack
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/word_access_start/$entry
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/word_access_start/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/word_access_start/word_0/rr
      -- 
    rr_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(162), ack => ptr_deref_713_store_0_req_0); -- 
    testConfigure_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(129) & testConfigure_CP_0_elements(133) & testConfigure_CP_0_elements(137) & testConfigure_CP_0_elements(141) & testConfigure_CP_0_elements(145) & testConfigure_CP_0_elements(149) & testConfigure_CP_0_elements(153) & testConfigure_CP_0_elements(157) & testConfigure_CP_0_elements(161);
      gj_testConfigure_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/word_access_start/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/word_access_start/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Sample/word_access_start/word_0/ra
      -- 
    ra_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_713_store_0_ack_0, ack => testConfigure_CP_0_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	295 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Update/word_access_complete/$exit
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Update/word_access_complete/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Update/word_access_complete/word_0/ca
      -- 
    ca_1930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_713_store_0_ack_1, ack => testConfigure_CP_0_elements(164)); -- 
    -- CP-element group 165:  branch  join  transition  place  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	126 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (10) 
      -- CP-element group 165: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726__exit__
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_727__entry__
      -- CP-element group 165: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_727_dead_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_727_eval_test/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_727_eval_test/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_727_eval_test/branch_req
      -- CP-element group 165: 	 branch_block_stmt_33/R_exitcond10_728_place
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_727_if_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_727_else_link/$entry
      -- 
    branch_req_1938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(165), ack => if_stmt_727_branch_req_0); -- 
    testConfigure_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(126) & testConfigure_CP_0_elements(164);
      gj_testConfigure_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  merge  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	289 
    -- CP-element group 166:  members (13) 
      -- CP-element group 166: 	 branch_block_stmt_33/merge_stmt_507__exit__
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader
      -- CP-element group 166: 	 branch_block_stmt_33/if_stmt_727_if_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_33/if_stmt_727_if_link/if_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 166: 	 branch_block_stmt_33/merge_stmt_507_PhiReqMerge
      -- CP-element group 166: 	 branch_block_stmt_33/merge_stmt_507_PhiAck/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/merge_stmt_507_PhiAck/$exit
      -- CP-element group 166: 	 branch_block_stmt_33/merge_stmt_507_PhiAck/dummy
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_727_branch_ack_1, ack => testConfigure_CP_0_elements(166)); -- 
    -- CP-element group 167:  fork  transition  place  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	291 
    -- CP-element group 167: 	292 
    -- CP-element group 167:  members (12) 
      -- CP-element group 167: 	 branch_block_stmt_33/if_stmt_727_else_link/$exit
      -- CP-element group 167: 	 branch_block_stmt_33/if_stmt_727_else_link/else_choice_transition
      -- CP-element group 167: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67
      -- CP-element group 167: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/$entry
      -- CP-element group 167: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/$entry
      -- CP-element group 167: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/$entry
      -- CP-element group 167: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/$entry
      -- CP-element group 167: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/SplitProtocol/$entry
      -- CP-element group 167: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/SplitProtocol/Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/SplitProtocol/Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/SplitProtocol/Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_727_branch_ack_0, ack => testConfigure_CP_0_elements(167)); -- 
    rr_3091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => type_cast_570_inst_req_0); -- 
    cr_3096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => type_cast_570_inst_req_1); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	123 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_Sample/ra
      -- 
    ra_1961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_0, ack => testConfigure_CP_0_elements(168)); -- 
    -- CP-element group 169:  transition  place  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	123 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	296 
    -- CP-element group 169:  members (9) 
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771__exit__
      -- CP-element group 169: 	 branch_block_stmt_33/bbx_xnph210_forx_xbody126
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/$exit
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_738_to_assign_stmt_771/type_cast_751_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_33/bbx_xnph210_forx_xbody126_PhiReq/$entry
      -- CP-element group 169: 	 branch_block_stmt_33/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_774/$entry
      -- CP-element group 169: 	 branch_block_stmt_33/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/$entry
      -- 
    ca_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_1, ack => testConfigure_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	301 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	209 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_final_index_sum_regn_sample_complete
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_final_index_sum_regn_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_final_index_sum_regn_Sample/ack
      -- 
    ack_1995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_786_index_offset_ack_0, ack => testConfigure_CP_0_elements(170)); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	301 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (11) 
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_root_address_calculated
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_offset_calculated
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_final_index_sum_regn_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_final_index_sum_regn_Update/ack
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_base_plus_offset/$entry
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_base_plus_offset/$exit
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_base_plus_offset/sum_rename_req
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_base_plus_offset/sum_rename_ack
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_request/$entry
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_request/req
      -- 
    ack_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_786_index_offset_ack_1, ack => testConfigure_CP_0_elements(171)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(171), ack => addr_of_787_final_reg_req_0); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_request/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_request/ack
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_787_final_reg_ack_0, ack => testConfigure_CP_0_elements(172)); -- 
    -- CP-element group 173:  fork  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	301 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	206 
    -- CP-element group 173:  members (19) 
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_word_addrgen/root_register_ack
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_word_addrgen/root_register_req
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_word_addrgen/$exit
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_word_addrgen/$entry
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_base_plus_offset/sum_rename_ack
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_base_plus_offset/sum_rename_req
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_base_plus_offset/$exit
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_base_plus_offset/$entry
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_base_addr_resize/base_resize_ack
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_base_addr_resize/base_resize_req
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_base_addr_resize/$exit
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_base_addr_resize/$entry
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_base_address_resized
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_root_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_word_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_base_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_complete/$exit
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_complete/ack
      -- 
    ack_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_787_final_reg_ack_1, ack => testConfigure_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	301 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (6) 
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_update_start_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_Sample/ra
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_Update/cr
      -- 
    ra_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_790_inst_ack_0, ack => testConfigure_CP_0_elements(174)); -- 
    cr_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(174), ack => RPIPE_ConvTranspose_input_pipe_790_inst_req_1); -- 
    -- CP-element group 175:  fork  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: 	178 
    -- CP-element group 175:  members (9) 
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_Update/ca
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_Sample/rr
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_Sample/rr
      -- 
    ca_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_790_inst_ack_1, ack => testConfigure_CP_0_elements(175)); -- 
    rr_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(175), ack => type_cast_794_inst_req_0); -- 
    rr_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(175), ack => RPIPE_ConvTranspose_input_pipe_803_inst_req_0); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_Sample/ra
      -- 
    ra_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_794_inst_ack_0, ack => testConfigure_CP_0_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	301 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	206 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_Update/ca
      -- 
    ca_2043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_794_inst_ack_1, ack => testConfigure_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	175 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (6) 
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_update_start_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_Sample/ra
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_Update/cr
      -- 
    ra_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_803_inst_ack_0, ack => testConfigure_CP_0_elements(178)); -- 
    cr_2056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(178), ack => RPIPE_ConvTranspose_input_pipe_803_inst_req_1); -- 
    -- CP-element group 179:  fork  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: 	182 
    -- CP-element group 179:  members (9) 
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_803_Update/ca
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_Sample/rr
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_Sample/rr
      -- 
    ca_2057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_803_inst_ack_1, ack => testConfigure_CP_0_elements(179)); -- 
    rr_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => type_cast_807_inst_req_0); -- 
    rr_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => RPIPE_ConvTranspose_input_pipe_821_inst_req_0); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_Sample/ra
      -- 
    ra_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_0, ack => testConfigure_CP_0_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	301 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	206 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_Update/ca
      -- 
    ca_2071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_1, ack => testConfigure_CP_0_elements(181)); -- 
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	179 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (6) 
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_update_start_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_Sample/ra
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_Update/cr
      -- 
    ra_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_821_inst_ack_0, ack => testConfigure_CP_0_elements(182)); -- 
    cr_2084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(182), ack => RPIPE_ConvTranspose_input_pipe_821_inst_req_1); -- 
    -- CP-element group 183:  fork  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183: 	186 
    -- CP-element group 183:  members (9) 
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_821_Update/ca
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_Sample/rr
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_Sample/rr
      -- 
    ca_2085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_821_inst_ack_1, ack => testConfigure_CP_0_elements(183)); -- 
    rr_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => type_cast_825_inst_req_0); -- 
    rr_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => RPIPE_ConvTranspose_input_pipe_839_inst_req_0); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_Sample/ra
      -- 
    ra_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_825_inst_ack_0, ack => testConfigure_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	301 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	206 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_Update/ca
      -- 
    ca_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_825_inst_ack_1, ack => testConfigure_CP_0_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	183 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_update_start_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_Sample/ra
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_Update/cr
      -- 
    ra_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_839_inst_ack_0, ack => testConfigure_CP_0_elements(186)); -- 
    cr_2112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(186), ack => RPIPE_ConvTranspose_input_pipe_839_inst_req_1); -- 
    -- CP-element group 187:  fork  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: 	190 
    -- CP-element group 187:  members (9) 
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_839_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_Sample/rr
      -- 
    ca_2113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_839_inst_ack_1, ack => testConfigure_CP_0_elements(187)); -- 
    rr_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => type_cast_843_inst_req_0); -- 
    rr_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => RPIPE_ConvTranspose_input_pipe_857_inst_req_0); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_Sample/ra
      -- 
    ra_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_0, ack => testConfigure_CP_0_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	301 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	206 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_Update/ca
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_update_completed_
      -- 
    ca_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_1, ack => testConfigure_CP_0_elements(189)); -- 
    -- CP-element group 190:  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	187 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (6) 
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_Sample/ra
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_update_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_Sample/$exit
      -- 
    ra_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_857_inst_ack_0, ack => testConfigure_CP_0_elements(190)); -- 
    cr_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(190), ack => RPIPE_ConvTranspose_input_pipe_857_inst_req_1); -- 
    -- CP-element group 191:  fork  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191: 	194 
    -- CP-element group 191:  members (9) 
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_Update/ca
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_Sample/rr
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_857_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_Sample/rr
      -- 
    ca_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_857_inst_ack_1, ack => testConfigure_CP_0_elements(191)); -- 
    rr_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => type_cast_861_inst_req_0); -- 
    rr_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => RPIPE_ConvTranspose_input_pipe_875_inst_req_0); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_Sample/ra
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_Sample/$exit
      -- 
    ra_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_861_inst_ack_0, ack => testConfigure_CP_0_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	301 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	206 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_Update/ca
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_update_completed_
      -- 
    ca_2155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_861_inst_ack_1, ack => testConfigure_CP_0_elements(193)); -- 
    -- CP-element group 194:  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	191 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_update_start_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_Update/cr
      -- 
    ra_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_875_inst_ack_0, ack => testConfigure_CP_0_elements(194)); -- 
    cr_2168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(194), ack => RPIPE_ConvTranspose_input_pipe_875_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195: 	198 
    -- CP-element group 195:  members (9) 
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_875_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_Sample/rr
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_Sample/rr
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_sample_start_
      -- 
    ca_2169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_875_inst_ack_1, ack => testConfigure_CP_0_elements(195)); -- 
    rr_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => type_cast_879_inst_req_0); -- 
    rr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => RPIPE_ConvTranspose_input_pipe_893_inst_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_Sample/ra
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_sample_completed_
      -- 
    ra_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_879_inst_ack_0, ack => testConfigure_CP_0_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	301 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	206 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_Update/ca
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_update_completed_
      -- 
    ca_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_879_inst_ack_1, ack => testConfigure_CP_0_elements(197)); -- 
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	195 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_Update/cr
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_update_start_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_sample_completed_
      -- 
    ra_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_893_inst_ack_0, ack => testConfigure_CP_0_elements(198)); -- 
    cr_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(198), ack => RPIPE_ConvTranspose_input_pipe_893_inst_req_1); -- 
    -- CP-element group 199:  fork  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: 	202 
    -- CP-element group 199:  members (9) 
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_Update/ca
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_893_update_completed_
      -- 
    ca_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_893_inst_ack_1, ack => testConfigure_CP_0_elements(199)); -- 
    rr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => type_cast_897_inst_req_0); -- 
    rr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => RPIPE_ConvTranspose_input_pipe_911_inst_req_0); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_sample_completed_
      -- 
    ra_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_897_inst_ack_0, ack => testConfigure_CP_0_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	301 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	206 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_Update/ca
      -- 
    ca_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_897_inst_ack_1, ack => testConfigure_CP_0_elements(201)); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	199 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_sample_completed_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_update_start_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_Sample/ra
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_Update/cr
      -- 
    ra_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_911_inst_ack_0, ack => testConfigure_CP_0_elements(202)); -- 
    cr_2224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(202), ack => RPIPE_ConvTranspose_input_pipe_911_inst_req_1); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_Sample/rr
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_911_Update/ca
      -- 
    ca_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_911_inst_ack_1, ack => testConfigure_CP_0_elements(203)); -- 
    rr_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(203), ack => type_cast_915_inst_req_0); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_Sample/ra
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_sample_completed_
      -- 
    ra_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_915_inst_ack_0, ack => testConfigure_CP_0_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	301 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_Update/ca
      -- 
    ca_2239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_915_inst_ack_1, ack => testConfigure_CP_0_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	173 
    -- CP-element group 206: 	177 
    -- CP-element group 206: 	181 
    -- CP-element group 206: 	185 
    -- CP-element group 206: 	189 
    -- CP-element group 206: 	193 
    -- CP-element group 206: 	197 
    -- CP-element group 206: 	201 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (9) 
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/word_access_start/word_0/rr
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/word_access_start/word_0/$entry
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/word_access_start/$entry
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/ptr_deref_923_Split/split_ack
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/ptr_deref_923_Split/split_req
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/ptr_deref_923_Split/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/ptr_deref_923_Split/$entry
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/$entry
      -- 
    rr_2277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(206), ack => ptr_deref_923_store_0_req_0); -- 
    testConfigure_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(173) & testConfigure_CP_0_elements(177) & testConfigure_CP_0_elements(181) & testConfigure_CP_0_elements(185) & testConfigure_CP_0_elements(189) & testConfigure_CP_0_elements(193) & testConfigure_CP_0_elements(197) & testConfigure_CP_0_elements(201) & testConfigure_CP_0_elements(205);
      gj_testConfigure_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/word_access_start/word_0/ra
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/word_access_start/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/word_access_start/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Sample/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_sample_completed_
      -- 
    ra_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_923_store_0_ack_0, ack => testConfigure_CP_0_elements(207)); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	301 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Update/word_access_complete/word_0/ca
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Update/word_access_complete/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Update/word_access_complete/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_update_completed_
      -- 
    ca_2289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_923_store_0_ack_1, ack => testConfigure_CP_0_elements(208)); -- 
    -- CP-element group 209:  branch  join  transition  place  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	170 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (10) 
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_937_else_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936__exit__
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_937__entry__
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_937_if_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_937_eval_test/branch_req
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_937_eval_test/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_937_eval_test/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_937_dead_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/R_exitcond19_938_place
      -- CP-element group 209: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/$exit
      -- 
    branch_req_2297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(209), ack => if_stmt_937_branch_req_0); -- 
    testConfigure_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(170) & testConfigure_CP_0_elements(208);
      gj_testConfigure_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  merge  transition  place  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	302 
    -- CP-element group 210:  members (13) 
      -- CP-element group 210: 	 branch_block_stmt_33/if_stmt_937_if_link/if_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_33/merge_stmt_943__exit__
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xend180x_xloopexit_forx_xend180
      -- CP-element group 210: 	 branch_block_stmt_33/if_stmt_937_if_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody126_forx_xend180x_xloopexit
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody126_forx_xend180x_xloopexit_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody126_forx_xend180x_xloopexit_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_33/merge_stmt_943_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_33/merge_stmt_943_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/merge_stmt_943_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_33/merge_stmt_943_PhiAck/dummy
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xend180x_xloopexit_forx_xend180_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xend180x_xloopexit_forx_xend180_PhiReq/$exit
      -- 
    if_choice_transition_2302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_937_branch_ack_1, ack => testConfigure_CP_0_elements(210)); -- 
    -- CP-element group 211:  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	297 
    -- CP-element group 211: 	298 
    -- CP-element group 211:  members (12) 
      -- CP-element group 211: 	 branch_block_stmt_33/if_stmt_937_else_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_33/if_stmt_937_else_link/else_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126
      -- CP-element group 211: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/$entry
      -- CP-element group 211: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/$entry
      -- CP-element group 211: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/$entry
      -- CP-element group 211: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/SplitProtocol/$entry
      -- CP-element group 211: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/SplitProtocol/Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/SplitProtocol/Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/SplitProtocol/Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_937_branch_ack_0, ack => testConfigure_CP_0_elements(211)); -- 
    rr_3145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => type_cast_780_inst_req_0); -- 
    cr_3150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => type_cast_780_inst_req_1); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	303 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (5) 
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Sample/word_access_start/$exit
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Sample/word_access_start/word_0/$exit
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Sample/word_access_start/word_0/ra
      -- 
    ra_2345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_956_load_0_ack_0, ack => testConfigure_CP_0_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	303 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	218 
    -- CP-element group 213:  members (9) 
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/word_access_complete/$exit
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/ptr_deref_956_Merge/merge_ack
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/ptr_deref_956_Merge/merge_req
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/ptr_deref_956_Merge/$exit
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/ptr_deref_956_Merge/$entry
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/word_access_complete/word_0/ca
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/word_access_complete/word_0/$exit
      -- 
    ca_2356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_956_load_0_ack_1, ack => testConfigure_CP_0_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	303 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (5) 
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_sample_completed_
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Sample/word_access_start/word_0/ra
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Sample/word_access_start/word_0/$exit
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Sample/word_access_start/$exit
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Sample/$exit
      -- 
    ra_2395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_968_load_0_ack_0, ack => testConfigure_CP_0_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	303 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	218 
    -- CP-element group 215:  members (9) 
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/ptr_deref_968_Merge/merge_ack
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/ptr_deref_968_Merge/merge_req
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/ptr_deref_968_Merge/$exit
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/ptr_deref_968_Merge/$entry
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/word_access_complete/word_0/ca
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/word_access_complete/word_0/$exit
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/word_access_complete/$exit
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/$exit
      -- 
    ca_2406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_968_load_0_ack_1, ack => testConfigure_CP_0_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	303 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (5) 
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Sample/word_access_start/$exit
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Sample/word_access_start/word_0/$exit
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Sample/word_access_start/word_0/ra
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_sample_completed_
      -- 
    ra_2445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_980_load_0_ack_0, ack => testConfigure_CP_0_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	303 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (9) 
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/ptr_deref_980_Merge/merge_ack
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/ptr_deref_980_Merge/merge_req
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/ptr_deref_980_Merge/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/ptr_deref_980_Merge/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/word_access_complete/word_0/ca
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/word_access_complete/word_0/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/word_access_complete/$exit
      -- 
    ca_2456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_980_load_0_ack_1, ack => testConfigure_CP_0_elements(217)); -- 
    -- CP-element group 218:  branch  join  transition  place  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	213 
    -- CP-element group 218: 	215 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (10) 
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997__exit__
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_998__entry__
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_998_eval_test/branch_req
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_998_eval_test/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/R_cmp191204_999_place
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_998_eval_test/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_998_if_link/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_998_else_link/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_998_dead_link/$entry
      -- 
    branch_req_2469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(218), ack => if_stmt_998_branch_req_0); -- 
    testConfigure_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(213) & testConfigure_CP_0_elements(215) & testConfigure_CP_0_elements(217);
      gj_testConfigure_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219: 	222 
    -- CP-element group 219:  members (18) 
      -- CP-element group 219: 	 branch_block_stmt_33/merge_stmt_1004__exit__
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039__entry__
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_update_start_
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_Sample/rr
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_Update/cr
      -- CP-element group 219: 	 branch_block_stmt_33/if_stmt_998_if_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_33/if_stmt_998_if_link/if_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/$entry
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend180_bbx_xnph
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend180_bbx_xnph_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend180_bbx_xnph_PhiReq/$exit
      -- CP-element group 219: 	 branch_block_stmt_33/merge_stmt_1004_PhiReqMerge
      -- CP-element group 219: 	 branch_block_stmt_33/merge_stmt_1004_PhiAck/$entry
      -- CP-element group 219: 	 branch_block_stmt_33/merge_stmt_1004_PhiAck/$exit
      -- CP-element group 219: 	 branch_block_stmt_33/merge_stmt_1004_PhiAck/dummy
      -- 
    if_choice_transition_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_998_branch_ack_1, ack => testConfigure_CP_0_elements(219)); -- 
    rr_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => type_cast_1025_inst_req_0); -- 
    cr_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => type_cast_1025_inst_req_1); -- 
    -- CP-element group 220:  transition  place  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	310 
    -- CP-element group 220:  members (5) 
      -- CP-element group 220: 	 branch_block_stmt_33/forx_xend180_forx_xend200
      -- CP-element group 220: 	 branch_block_stmt_33/if_stmt_998_else_link/else_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_33/if_stmt_998_else_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_33/forx_xend180_forx_xend200_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_33/forx_xend180_forx_xend200_PhiReq/$exit
      -- 
    else_choice_transition_2478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_998_branch_ack_0, ack => testConfigure_CP_0_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_Sample/ra
      -- 
    ra_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_0, ack => testConfigure_CP_0_elements(221)); -- 
    -- CP-element group 222:  transition  place  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	219 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	304 
    -- CP-element group 222:  members (9) 
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039__exit__
      -- CP-element group 222: 	 branch_block_stmt_33/bbx_xnph_forx_xbody193
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/type_cast_1025_Update/ca
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_1010_to_assign_stmt_1039/$exit
      -- CP-element group 222: 	 branch_block_stmt_33/bbx_xnph_forx_xbody193_PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_33/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1042/$entry
      -- CP-element group 222: 	 branch_block_stmt_33/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/$entry
      -- 
    ca_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_1, ack => testConfigure_CP_0_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	309 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	229 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_final_index_sum_regn_Sample/ack
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_final_index_sum_regn_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_final_index_sum_regn_sample_complete
      -- 
    ack_2526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1054_index_offset_ack_0, ack => testConfigure_CP_0_elements(223)); -- 
    -- CP-element group 224:  transition  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	309 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (11) 
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_base_plus_offset/sum_rename_ack
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_base_plus_offset/sum_rename_req
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_request/$entry
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_sample_start_
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_request/req
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_base_plus_offset/$exit
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_base_plus_offset/$entry
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_final_index_sum_regn_Update/ack
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_final_index_sum_regn_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_offset_calculated
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_root_address_calculated
      -- 
    ack_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1054_index_offset_ack_1, ack => testConfigure_CP_0_elements(224)); -- 
    req_2540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(224), ack => addr_of_1055_final_reg_req_0); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_request/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_request/ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_sample_completed_
      -- 
    ack_2541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1055_final_reg_ack_0, ack => testConfigure_CP_0_elements(225)); -- 
    -- CP-element group 226:  join  fork  transition  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	309 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (28) 
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_base_addr_resize/base_resize_req
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_word_addrgen/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_base_addr_resize/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_word_addrgen/$entry
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_base_plus_offset/sum_rename_ack
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_base_addr_resize/$entry
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/word_access_start/word_0/$entry
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_base_address_resized
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_base_plus_offset/sum_rename_req
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_base_plus_offset/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/word_access_start/$entry
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_root_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_base_plus_offset/$entry
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/ptr_deref_1058_Split/split_ack
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_word_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/ptr_deref_1058_Split/split_req
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_word_addrgen/root_register_ack
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/ptr_deref_1058_Split/$entry
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/ptr_deref_1058_Split/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_complete/ack
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_base_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_word_addrgen/root_register_req
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_complete/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_base_addr_resize/base_resize_ack
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/word_access_start/word_0/rr
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_update_completed_
      -- 
    ack_2546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1055_final_reg_ack_1, ack => testConfigure_CP_0_elements(226)); -- 
    rr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(226), ack => ptr_deref_1058_store_0_req_0); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/word_access_start/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/word_access_start/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Sample/word_access_start/word_0/ra
      -- 
    ra_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1058_store_0_ack_0, ack => testConfigure_CP_0_elements(227)); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	309 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Update/word_access_complete/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Update/word_access_complete/word_0/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Update/word_access_complete/word_0/ca
      -- 
    ca_2596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1058_store_0_ack_1, ack => testConfigure_CP_0_elements(228)); -- 
    -- CP-element group 229:  branch  join  transition  place  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	223 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (10) 
      -- CP-element group 229: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072__exit__
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_1073__entry__
      -- CP-element group 229: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_1073_dead_link/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_1073_eval_test/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_1073_eval_test/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_1073_eval_test/branch_req
      -- CP-element group 229: 	 branch_block_stmt_33/R_exitcond20_1074_place
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_1073_if_link/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_1073_else_link/$entry
      -- 
    branch_req_2604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => if_stmt_1073_branch_req_0); -- 
    testConfigure_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(223) & testConfigure_CP_0_elements(228);
      gj_testConfigure_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  merge  transition  place  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	310 
    -- CP-element group 230:  members (13) 
      -- CP-element group 230: 	 branch_block_stmt_33/merge_stmt_1079__exit__
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xend200x_xloopexit_forx_xend200
      -- CP-element group 230: 	 branch_block_stmt_33/if_stmt_1073_if_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_33/if_stmt_1073_if_link/if_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody193_forx_xend200x_xloopexit
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody193_forx_xend200x_xloopexit_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody193_forx_xend200x_xloopexit_PhiReq/$exit
      -- CP-element group 230: 	 branch_block_stmt_33/merge_stmt_1079_PhiReqMerge
      -- CP-element group 230: 	 branch_block_stmt_33/merge_stmt_1079_PhiAck/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/merge_stmt_1079_PhiAck/$exit
      -- CP-element group 230: 	 branch_block_stmt_33/merge_stmt_1079_PhiAck/dummy
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xend200x_xloopexit_forx_xend200_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xend200x_xloopexit_forx_xend200_PhiReq/$exit
      -- 
    if_choice_transition_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1073_branch_ack_1, ack => testConfigure_CP_0_elements(230)); -- 
    -- CP-element group 231:  fork  transition  place  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	305 
    -- CP-element group 231: 	306 
    -- CP-element group 231:  members (12) 
      -- CP-element group 231: 	 branch_block_stmt_33/if_stmt_1073_else_link/$exit
      -- CP-element group 231: 	 branch_block_stmt_33/if_stmt_1073_else_link/else_choice_transition
      -- CP-element group 231: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193
      -- CP-element group 231: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/$entry
      -- CP-element group 231: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/$entry
      -- CP-element group 231: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/$entry
      -- CP-element group 231: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/$entry
      -- CP-element group 231: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/SplitProtocol/$entry
      -- CP-element group 231: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/SplitProtocol/Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/SplitProtocol/Sample/rr
      -- CP-element group 231: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/SplitProtocol/Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1073_branch_ack_0, ack => testConfigure_CP_0_elements(231)); -- 
    rr_3222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(231), ack => type_cast_1048_inst_req_0); -- 
    cr_3227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(231), ack => type_cast_1048_inst_req_1); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	310 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_Sample/ra
      -- 
    ra_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1084_inst_ack_0, ack => testConfigure_CP_0_elements(232)); -- 
    -- CP-element group 233:  transition  place  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	310 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (16) 
      -- CP-element group 233: 	 $exit
      -- CP-element group 233: 	 branch_block_stmt_33/$exit
      -- CP-element group 233: 	 branch_block_stmt_33/branch_block_stmt_33__exit__
      -- CP-element group 233: 	 branch_block_stmt_33/assign_stmt_1085__exit__
      -- CP-element group 233: 	 branch_block_stmt_33/return__
      -- CP-element group 233: 	 branch_block_stmt_33/merge_stmt_1087__exit__
      -- CP-element group 233: 	 branch_block_stmt_33/assign_stmt_1085/$exit
      -- CP-element group 233: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_Update/ca
      -- CP-element group 233: 	 branch_block_stmt_33/return___PhiReq/$entry
      -- CP-element group 233: 	 branch_block_stmt_33/return___PhiReq/$exit
      -- CP-element group 233: 	 branch_block_stmt_33/merge_stmt_1087_PhiReqMerge
      -- CP-element group 233: 	 branch_block_stmt_33/merge_stmt_1087_PhiAck/$entry
      -- CP-element group 233: 	 branch_block_stmt_33/merge_stmt_1087_PhiAck/$exit
      -- CP-element group 233: 	 branch_block_stmt_33/merge_stmt_1087_PhiAck/dummy
      -- 
    ca_2632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1084_inst_ack_1, ack => testConfigure_CP_0_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	32 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (2) 
      -- CP-element group 234: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/SplitProtocol/Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/SplitProtocol/Sample/ra
      -- 
    ra_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_0, ack => testConfigure_CP_0_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	32 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/SplitProtocol/Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/SplitProtocol/Update/ca
      -- 
    ca_2669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_1, ack => testConfigure_CP_0_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	240 
    -- CP-element group 236:  members (5) 
      -- CP-element group 236: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/$exit
      -- CP-element group 236: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/$exit
      -- CP-element group 236: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/$exit
      -- CP-element group 236: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_77/SplitProtocol/$exit
      -- CP-element group 236: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_req
      -- 
    phi_stmt_74_req_2670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_74_req_2670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(236), ack => phi_stmt_74_req_0); -- 
    testConfigure_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(234) & testConfigure_CP_0_elements(235);
      gj_testConfigure_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	32 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (2) 
      -- CP-element group 237: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/SplitProtocol/Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/SplitProtocol/Sample/ra
      -- 
    ra_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_84_inst_ack_0, ack => testConfigure_CP_0_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	32 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (2) 
      -- CP-element group 238: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/SplitProtocol/Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/SplitProtocol/Update/ca
      -- 
    ca_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_84_inst_ack_1, ack => testConfigure_CP_0_elements(238)); -- 
    -- CP-element group 239:  join  transition  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (5) 
      -- CP-element group 239: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/$exit
      -- CP-element group 239: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/$exit
      -- CP-element group 239: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/$exit
      -- CP-element group 239: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_84/SplitProtocol/$exit
      -- CP-element group 239: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_req
      -- 
    phi_stmt_81_req_2693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_81_req_2693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(239), ack => phi_stmt_81_req_0); -- 
    testConfigure_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(237) & testConfigure_CP_0_elements(238);
      gj_testConfigure_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  join  transition  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	236 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	246 
    -- CP-element group 240:  members (1) 
      -- CP-element group 240: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(236) & testConfigure_CP_0_elements(239);
      gj_testConfigure_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  transition  output  delay-element  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	14 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	245 
    -- CP-element group 241:  members (4) 
      -- CP-element group 241: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_74/$exit
      -- CP-element group 241: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/$exit
      -- CP-element group 241: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_sources/type_cast_80_konst_delay_trans
      -- CP-element group 241: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_74/phi_stmt_74_req
      -- 
    phi_stmt_74_req_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_74_req_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => phi_stmt_74_req_1); -- 
    -- Element group testConfigure_CP_0_elements(241) is a control-delay.
    cp_element_241_delay: control_delay_element  generic map(name => " 241_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(14), ack => testConfigure_CP_0_elements(241), clk => clk, reset =>reset);
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	14 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/SplitProtocol/Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/SplitProtocol/Sample/ra
      -- 
    ra_2721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_86_inst_ack_0, ack => testConfigure_CP_0_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	14 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/SplitProtocol/Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/SplitProtocol/Update/ca
      -- 
    ca_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_86_inst_ack_1, ack => testConfigure_CP_0_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (5) 
      -- CP-element group 244: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/$exit
      -- CP-element group 244: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/$exit
      -- CP-element group 244: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/$exit
      -- CP-element group 244: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_sources/type_cast_86/SplitProtocol/$exit
      -- CP-element group 244: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_81/phi_stmt_81_req
      -- 
    phi_stmt_81_req_2727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_81_req_2727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => phi_stmt_81_req_1); -- 
    testConfigure_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(242) & testConfigure_CP_0_elements(243);
      gj_testConfigure_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	241 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (1) 
      -- CP-element group 245: 	 branch_block_stmt_33/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(241) & testConfigure_CP_0_elements(244);
      gj_testConfigure_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  merge  fork  transition  place  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	240 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (2) 
      -- CP-element group 246: 	 branch_block_stmt_33/merge_stmt_73_PhiReqMerge
      -- CP-element group 246: 	 branch_block_stmt_33/merge_stmt_73_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(246) <= OrReduce(testConfigure_CP_0_elements(240) & testConfigure_CP_0_elements(245));
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	249 
    -- CP-element group 247:  members (1) 
      -- CP-element group 247: 	 branch_block_stmt_33/merge_stmt_73_PhiAck/phi_stmt_74_ack
      -- 
    phi_stmt_74_ack_2732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_74_ack_0, ack => testConfigure_CP_0_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (1) 
      -- CP-element group 248: 	 branch_block_stmt_33/merge_stmt_73_PhiAck/phi_stmt_81_ack
      -- 
    phi_stmt_81_ack_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_81_ack_0, ack => testConfigure_CP_0_elements(248)); -- 
    -- CP-element group 249:  join  fork  transition  place  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	15 
    -- CP-element group 249: 	16 
    -- CP-element group 249: 	17 
    -- CP-element group 249: 	18 
    -- CP-element group 249: 	20 
    -- CP-element group 249: 	22 
    -- CP-element group 249: 	23 
    -- CP-element group 249: 	25 
    -- CP-element group 249: 	26 
    -- CP-element group 249: 	29 
    -- CP-element group 249:  members (61) 
      -- CP-element group 249: 	 branch_block_stmt_33/merge_stmt_73__exit__
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136__entry__
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_update_start_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_base_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_word_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_root_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_base_address_resized
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_base_addr_resize/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_base_addr_resize/$exit
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_update_start_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_96_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_update_start_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_resized_1
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_scaled_1
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_computed_1
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_resize_1/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_resize_1/$exit
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_resize_1/index_resize_req
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_resize_1/index_resize_ack
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_scale_1/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_scale_1/$exit
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_scale_1/scale_rename_req
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_index_scale_1/scale_rename_ack
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_final_index_sum_regn_update_start
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_final_index_sum_regn_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_final_index_sum_regn_Sample/req
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_final_index_sum_regn_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/array_obj_ref_102_final_index_sum_regn_Update/req
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/addr_of_103_complete/req
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_update_start_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Update/word_access_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Update/word_access_complete/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_106_Update/word_access_complete/word_0/cr
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_base_addr_resize/base_resize_req
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_base_addr_resize/base_resize_ack
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_base_plus_offset/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_base_plus_offset/$exit
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_base_plus_offset/sum_rename_req
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_base_plus_offset/sum_rename_ack
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_word_addrgen/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_word_addrgen/$exit
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_word_addrgen/root_register_req
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_word_addrgen/root_register_ack
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/word_access_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/word_access_complete/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/ptr_deref_123_Update/word_access_complete/word_0/cr
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/RPIPE_ConvTranspose_input_pipe_131_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_update_start_
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/assign_stmt_93_to_assign_stmt_136/type_cast_135_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_33/merge_stmt_73_PhiAck/$exit
      -- 
    rr_246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => type_cast_96_inst_req_0); -- 
    cr_251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => type_cast_96_inst_req_1); -- 
    req_277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => array_obj_ref_102_index_offset_req_0); -- 
    req_282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => array_obj_ref_102_index_offset_req_1); -- 
    req_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => addr_of_103_final_reg_req_1); -- 
    cr_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => ptr_deref_106_store_0_req_1); -- 
    cr_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => ptr_deref_123_load_0_req_1); -- 
    rr_406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => RPIPE_ConvTranspose_input_pipe_131_inst_req_0); -- 
    cr_425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => type_cast_135_inst_req_1); -- 
    testConfigure_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(247) & testConfigure_CP_0_elements(248);
      gj_testConfigure_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	33 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/SplitProtocol/Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/SplitProtocol/Sample/ra
      -- 
    ra_2757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_147_inst_ack_0, ack => testConfigure_CP_0_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	33 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (2) 
      -- CP-element group 251: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/SplitProtocol/Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/SplitProtocol/Update/ca
      -- 
    ca_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_147_inst_ack_1, ack => testConfigure_CP_0_elements(251)); -- 
    -- CP-element group 252:  join  transition  place  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (8) 
      -- CP-element group 252: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 252: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/$exit
      -- CP-element group 252: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/$exit
      -- CP-element group 252: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/$exit
      -- CP-element group 252: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_sources/type_cast_147/SplitProtocol/$exit
      -- CP-element group 252: 	 branch_block_stmt_33/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_144/phi_stmt_144_req
      -- CP-element group 252: 	 branch_block_stmt_33/merge_stmt_143_PhiReqMerge
      -- CP-element group 252: 	 branch_block_stmt_33/merge_stmt_143_PhiAck/$entry
      -- 
    phi_stmt_144_req_2763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_144_req_2763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(252), ack => phi_stmt_144_req_0); -- 
    testConfigure_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(250) & testConfigure_CP_0_elements(251);
      gj_testConfigure_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	257 
    -- CP-element group 253: 	258 
    -- CP-element group 253:  members (13) 
      -- CP-element group 253: 	 branch_block_stmt_33/merge_stmt_143__exit__
      -- CP-element group 253: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend
      -- CP-element group 253: 	 branch_block_stmt_33/merge_stmt_143_PhiAck/$exit
      -- CP-element group 253: 	 branch_block_stmt_33/merge_stmt_143_PhiAck/phi_stmt_144_ack
      -- CP-element group 253: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/SplitProtocol/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/SplitProtocol/Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/SplitProtocol/Sample/rr
      -- CP-element group 253: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/SplitProtocol/Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/SplitProtocol/Update/cr
      -- 
    phi_stmt_144_ack_2768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_144_ack_0, ack => testConfigure_CP_0_elements(253)); -- 
    rr_2813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(253), ack => type_cast_156_inst_req_0); -- 
    cr_2818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(253), ack => type_cast_156_inst_req_1); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	13 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (2) 
      -- CP-element group 254: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/SplitProtocol/Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/SplitProtocol/Sample/ra
      -- 
    ra_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_154_inst_ack_0, ack => testConfigure_CP_0_elements(254)); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	13 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (2) 
      -- CP-element group 255: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/SplitProtocol/Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/SplitProtocol/Update/ca
      -- 
    ca_2793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_154_inst_ack_1, ack => testConfigure_CP_0_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	260 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/$exit
      -- CP-element group 256: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/$exit
      -- CP-element group 256: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/$exit
      -- CP-element group 256: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/$exit
      -- CP-element group 256: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_154/SplitProtocol/$exit
      -- CP-element group 256: 	 branch_block_stmt_33/entry_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_req
      -- 
    phi_stmt_151_req_2794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_151_req_2794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(256), ack => phi_stmt_151_req_0); -- 
    testConfigure_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(254) & testConfigure_CP_0_elements(255);
      gj_testConfigure_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	253 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (2) 
      -- CP-element group 257: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/SplitProtocol/Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/SplitProtocol/Sample/ra
      -- 
    ra_2814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_156_inst_ack_0, ack => testConfigure_CP_0_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	253 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (2) 
      -- CP-element group 258: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/SplitProtocol/Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/SplitProtocol/Update/ca
      -- 
    ca_2819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_156_inst_ack_1, ack => testConfigure_CP_0_elements(258)); -- 
    -- CP-element group 259:  join  transition  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_sources/type_cast_156/SplitProtocol/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_151/phi_stmt_151_req
      -- 
    phi_stmt_151_req_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_151_req_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => phi_stmt_151_req_1); -- 
    testConfigure_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(257) & testConfigure_CP_0_elements(258);
      gj_testConfigure_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  merge  transition  place  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	256 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (2) 
      -- CP-element group 260: 	 branch_block_stmt_33/merge_stmt_150_PhiReqMerge
      -- CP-element group 260: 	 branch_block_stmt_33/merge_stmt_150_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(260) <= OrReduce(testConfigure_CP_0_elements(256) & testConfigure_CP_0_elements(259));
    -- CP-element group 261:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	34 
    -- CP-element group 261: 	35 
    -- CP-element group 261:  members (35) 
      -- CP-element group 261: 	 branch_block_stmt_33/merge_stmt_150__exit__
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173__entry__
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_update_start_
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_base_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_word_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_root_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_base_address_resized
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_base_addr_resize/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_base_addr_resize/$exit
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_base_addr_resize/base_resize_req
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_base_addr_resize/base_resize_ack
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_base_plus_offset/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_base_plus_offset/$exit
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_base_plus_offset/sum_rename_req
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_base_plus_offset/sum_rename_ack
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_word_addrgen/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_word_addrgen/$exit
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_word_addrgen/root_register_req
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_word_addrgen/root_register_ack
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/ptr_deref_165_Split/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/ptr_deref_165_Split/$exit
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/ptr_deref_165_Split/split_req
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/ptr_deref_165_Split/split_ack
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/word_access_start/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/word_access_start/word_0/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Sample/word_access_start/word_0/rr
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Update/word_access_complete/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Update/word_access_complete/word_0/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/assign_stmt_163_to_assign_stmt_173/ptr_deref_165_Update/word_access_complete/word_0/cr
      -- CP-element group 261: 	 branch_block_stmt_33/merge_stmt_150_PhiAck/$exit
      -- CP-element group 261: 	 branch_block_stmt_33/merge_stmt_150_PhiAck/phi_stmt_151_ack
      -- 
    phi_stmt_151_ack_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_151_ack_0, ack => testConfigure_CP_0_elements(261)); -- 
    rr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(261), ack => ptr_deref_165_store_0_req_0); -- 
    cr_498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(261), ack => ptr_deref_165_store_0_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	56 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (2) 
      -- CP-element group 262: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/SplitProtocol/Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/SplitProtocol/Sample/ra
      -- 
    ra_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_186_inst_ack_0, ack => testConfigure_CP_0_elements(262)); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	56 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (2) 
      -- CP-element group 263: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/SplitProtocol/Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/SplitProtocol/Update/ca
      -- 
    ca_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_186_inst_ack_1, ack => testConfigure_CP_0_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_186/SplitProtocol/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_req
      -- 
    phi_stmt_183_req_2863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_183_req_2863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(264), ack => phi_stmt_183_req_0); -- 
    testConfigure_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(262) & testConfigure_CP_0_elements(263);
      gj_testConfigure_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  transition  output  delay-element  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	37 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (5) 
      -- CP-element group 265: 	 branch_block_stmt_33/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/$exit
      -- CP-element group 265: 	 branch_block_stmt_33/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_183/$exit
      -- CP-element group 265: 	 branch_block_stmt_33/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/$exit
      -- CP-element group 265: 	 branch_block_stmt_33/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_sources/type_cast_189_konst_delay_trans
      -- CP-element group 265: 	 branch_block_stmt_33/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_183/phi_stmt_183_req
      -- 
    phi_stmt_183_req_2874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_183_req_2874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(265), ack => phi_stmt_183_req_1); -- 
    -- Element group testConfigure_CP_0_elements(265) is a control-delay.
    cp_element_265_delay: control_delay_element  generic map(name => " 265_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(37), ack => testConfigure_CP_0_elements(265), clk => clk, reset =>reset);
    -- CP-element group 266:  merge  transition  place  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (2) 
      -- CP-element group 266: 	 branch_block_stmt_33/merge_stmt_182_PhiReqMerge
      -- CP-element group 266: 	 branch_block_stmt_33/merge_stmt_182_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(266) <= OrReduce(testConfigure_CP_0_elements(264) & testConfigure_CP_0_elements(265));
    -- CP-element group 267:  fork  transition  place  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	44 
    -- CP-element group 267: 	47 
    -- CP-element group 267: 	43 
    -- CP-element group 267: 	50 
    -- CP-element group 267: 	51 
    -- CP-element group 267: 	38 
    -- CP-element group 267: 	39 
    -- CP-element group 267: 	40 
    -- CP-element group 267: 	41 
    -- CP-element group 267: 	53 
    -- CP-element group 267:  members (62) 
      -- CP-element group 267: 	 branch_block_stmt_33/merge_stmt_182__exit__
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239__entry__
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_update_start_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_199_Update/cr
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_update_start_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_resized_1
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_scaled_1
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_computed_1
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_resize_1/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_resize_1/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_resize_1/index_resize_req
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_resize_1/index_resize_ack
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_scale_1/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_scale_1/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_scale_1/scale_rename_req
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_index_scale_1/scale_rename_ack
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_final_index_sum_regn_update_start
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_final_index_sum_regn_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_final_index_sum_regn_Sample/req
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_final_index_sum_regn_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/array_obj_ref_205_final_index_sum_regn_Update/req
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_complete/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/addr_of_206_complete/req
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/RPIPE_ConvTranspose_input_pipe_209_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_update_start_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/type_cast_213_Update/cr
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_update_start_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Update/word_access_complete/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Update/word_access_complete/word_0/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_216_Update/word_access_complete/word_0/cr
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_update_start_
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_base_address_calculated
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_word_address_calculated
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_root_address_calculated
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_base_address_resized
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_base_addr_resize/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_base_addr_resize/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_base_addr_resize/base_resize_req
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_base_addr_resize/base_resize_ack
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_base_plus_offset/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_base_plus_offset/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_base_plus_offset/sum_rename_req
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_base_plus_offset/sum_rename_ack
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_word_addrgen/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_word_addrgen/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_word_addrgen/root_register_req
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_word_addrgen/root_register_ack
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/word_access_complete/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/word_access_complete/word_0/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/assign_stmt_196_to_assign_stmt_239/ptr_deref_233_Update/word_access_complete/word_0/cr
      -- CP-element group 267: 	 branch_block_stmt_33/merge_stmt_182_PhiAck/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/merge_stmt_182_PhiAck/phi_stmt_183_ack
      -- 
    phi_stmt_183_ack_2879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_183_ack_0, ack => testConfigure_CP_0_elements(267)); -- 
    rr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => type_cast_199_inst_req_0); -- 
    cr_534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => type_cast_199_inst_req_1); -- 
    req_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => array_obj_ref_205_index_offset_req_0); -- 
    req_565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => array_obj_ref_205_index_offset_req_1); -- 
    req_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => addr_of_206_final_reg_req_1); -- 
    rr_589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => RPIPE_ConvTranspose_input_pipe_209_inst_req_0); -- 
    cr_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => type_cast_213_inst_req_1); -- 
    cr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => ptr_deref_216_store_0_req_1); -- 
    cr_703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => ptr_deref_233_load_0_req_1); -- 
    -- CP-element group 268:  merge  fork  transition  place  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	36 
    -- CP-element group 268: 	57 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	58 
    -- CP-element group 268: 	61 
    -- CP-element group 268:  members (13) 
      -- CP-element group 268: 	 branch_block_stmt_33/merge_stmt_248__exit__
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255__entry__
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/$entry
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/RPIPE_ConvTranspose_input_pipe_250_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_update_start_
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_Update/$entry
      -- CP-element group 268: 	 branch_block_stmt_33/assign_stmt_251_to_assign_stmt_255/type_cast_254_Update/cr
      -- CP-element group 268: 	 branch_block_stmt_33/merge_stmt_248_PhiReqMerge
      -- CP-element group 268: 	 branch_block_stmt_33/merge_stmt_248_PhiAck/$entry
      -- CP-element group 268: 	 branch_block_stmt_33/merge_stmt_248_PhiAck/$exit
      -- CP-element group 268: 	 branch_block_stmt_33/merge_stmt_248_PhiAck/dummy
      -- 
    rr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(268), ack => RPIPE_ConvTranspose_input_pipe_250_inst_req_0); -- 
    cr_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(268), ack => type_cast_254_inst_req_1); -- 
    testConfigure_CP_0_elements(268) <= OrReduce(testConfigure_CP_0_elements(36) & testConfigure_CP_0_elements(57));
    -- CP-element group 269:  transition  output  delay-element  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	61 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	273 
    -- CP-element group 269:  members (4) 
      -- CP-element group 269: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_258/$exit
      -- CP-element group 269: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/$exit
      -- CP-element group 269: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_262_konst_delay_trans
      -- CP-element group 269: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_req
      -- 
    phi_stmt_258_req_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_258_req_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(269), ack => phi_stmt_258_req_0); -- 
    -- Element group testConfigure_CP_0_elements(269) is a control-delay.
    cp_element_269_delay: control_delay_element  generic map(name => " 269_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(61), ack => testConfigure_CP_0_elements(269), clk => clk, reset =>reset);
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	61 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (2) 
      -- CP-element group 270: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/SplitProtocol/Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/SplitProtocol/Sample/ra
      -- 
    ra_2930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_268_inst_ack_0, ack => testConfigure_CP_0_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	61 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (2) 
      -- CP-element group 271: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/SplitProtocol/Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/SplitProtocol/Update/ca
      -- 
    ca_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_268_inst_ack_1, ack => testConfigure_CP_0_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (5) 
      -- CP-element group 272: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/$exit
      -- CP-element group 272: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/$exit
      -- CP-element group 272: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/$exit
      -- CP-element group 272: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_268/SplitProtocol/$exit
      -- CP-element group 272: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_req
      -- 
    phi_stmt_265_req_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_265_req_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(272), ack => phi_stmt_265_req_0); -- 
    testConfigure_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(270) & testConfigure_CP_0_elements(271);
      gj_testConfigure_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	269 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	281 
    -- CP-element group 273:  members (1) 
      -- CP-element group 273: 	 branch_block_stmt_33/bbx_xnph221_forx_xbody28_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(269) & testConfigure_CP_0_elements(272);
      gj_testConfigure_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	72 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/SplitProtocol/Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/SplitProtocol/Sample/ra
      -- 
    ra_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_264_inst_ack_0, ack => testConfigure_CP_0_elements(274)); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	72 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (2) 
      -- CP-element group 275: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/SplitProtocol/Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/SplitProtocol/Update/ca
      -- 
    ca_2961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_264_inst_ack_1, ack => testConfigure_CP_0_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	280 
    -- CP-element group 276:  members (5) 
      -- CP-element group 276: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/$exit
      -- CP-element group 276: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/$exit
      -- CP-element group 276: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/$exit
      -- CP-element group 276: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_sources/type_cast_264/SplitProtocol/$exit
      -- CP-element group 276: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_258/phi_stmt_258_req
      -- 
    phi_stmt_258_req_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_258_req_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(276), ack => phi_stmt_258_req_1); -- 
    testConfigure_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(274) & testConfigure_CP_0_elements(275);
      gj_testConfigure_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	72 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (2) 
      -- CP-element group 277: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/SplitProtocol/Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/SplitProtocol/Sample/ra
      -- 
    ra_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_270_inst_ack_0, ack => testConfigure_CP_0_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	72 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (2) 
      -- CP-element group 278: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/SplitProtocol/Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/SplitProtocol/Update/ca
      -- 
    ca_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_270_inst_ack_1, ack => testConfigure_CP_0_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (5) 
      -- CP-element group 279: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/$exit
      -- CP-element group 279: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/$exit
      -- CP-element group 279: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/$exit
      -- CP-element group 279: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_sources/type_cast_270/SplitProtocol/$exit
      -- CP-element group 279: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_265/phi_stmt_265_req
      -- 
    phi_stmt_265_req_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_265_req_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => phi_stmt_265_req_1); -- 
    testConfigure_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(277) & testConfigure_CP_0_elements(278);
      gj_testConfigure_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  join  transition  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	276 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (1) 
      -- CP-element group 280: 	 branch_block_stmt_33/forx_xbody28_forx_xbody28_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(276) & testConfigure_CP_0_elements(279);
      gj_testConfigure_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  merge  fork  transition  place  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	273 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (2) 
      -- CP-element group 281: 	 branch_block_stmt_33/merge_stmt_257_PhiReqMerge
      -- CP-element group 281: 	 branch_block_stmt_33/merge_stmt_257_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(281) <= OrReduce(testConfigure_CP_0_elements(273) & testConfigure_CP_0_elements(280));
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_33/merge_stmt_257_PhiAck/phi_stmt_258_ack
      -- 
    phi_stmt_258_ack_2990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_258_ack_0, ack => testConfigure_CP_0_elements(282)); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (1) 
      -- CP-element group 283: 	 branch_block_stmt_33/merge_stmt_257_PhiAck/phi_stmt_265_ack
      -- 
    phi_stmt_265_ack_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_265_ack_0, ack => testConfigure_CP_0_elements(283)); -- 
    -- CP-element group 284:  join  fork  transition  place  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	62 
    -- CP-element group 284: 	63 
    -- CP-element group 284: 	65 
    -- CP-element group 284: 	66 
    -- CP-element group 284: 	69 
    -- CP-element group 284:  members (42) 
      -- CP-element group 284: 	 branch_block_stmt_33/merge_stmt_257__exit__
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299__entry__
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_base_plus_offset/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_base_plus_offset/$exit
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_base_plus_offset/sum_rename_req
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_base_plus_offset/sum_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_request/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_request/req
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_complete/req
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_update_start_
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/addr_of_275_update_start_
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_root_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_offset_calculated
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_resized_0
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_scaled_0
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_computed_0
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_resize_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_resize_0/$exit
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_resize_0/index_resize_req
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_resize_0/index_resize_ack
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_scale_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_scale_0/$exit
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_scale_0/scale_rename_req
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_index_scale_0/scale_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_final_index_sum_regn/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_final_index_sum_regn/$exit
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_final_index_sum_regn/req
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/array_obj_ref_274_final_index_sum_regn/ack
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Update/word_access_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Update/word_access_complete/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/ptr_deref_278_Update/word_access_complete/word_0/cr
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/RPIPE_ConvTranspose_input_pipe_282_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_update_start_
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/assign_stmt_276_to_assign_stmt_299/type_cast_286_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_33/merge_stmt_257_PhiAck/$exit
      -- 
    req_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => addr_of_275_final_reg_req_0); -- 
    req_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => addr_of_275_final_reg_req_1); -- 
    cr_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => ptr_deref_278_store_0_req_1); -- 
    rr_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => RPIPE_ConvTranspose_input_pipe_282_inst_req_0); -- 
    cr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => type_cast_286_inst_req_1); -- 
    testConfigure_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(282) & testConfigure_CP_0_elements(283);
      gj_testConfigure_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	71 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (2) 
      -- CP-element group 285: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/SplitProtocol/Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/SplitProtocol/Sample/ra
      -- 
    ra_3015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_310_inst_ack_0, ack => testConfigure_CP_0_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	71 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/SplitProtocol/Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/SplitProtocol/Update/ca
      -- 
    ca_3020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_310_inst_ack_1, ack => testConfigure_CP_0_elements(286)); -- 
    -- CP-element group 287:  join  transition  place  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (8) 
      -- CP-element group 287: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/$exit
      -- CP-element group 287: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/$exit
      -- CP-element group 287: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/$exit
      -- CP-element group 287: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/$exit
      -- CP-element group 287: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_sources/type_cast_310/SplitProtocol/$exit
      -- CP-element group 287: 	 branch_block_stmt_33/forx_xbody28_forx_xend37_PhiReq/phi_stmt_307/phi_stmt_307_req
      -- CP-element group 287: 	 branch_block_stmt_33/merge_stmt_306_PhiReqMerge
      -- CP-element group 287: 	 branch_block_stmt_33/merge_stmt_306_PhiAck/$entry
      -- 
    phi_stmt_307_req_3021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_307_req_3021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => phi_stmt_307_req_0); -- 
    testConfigure_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(285) & testConfigure_CP_0_elements(286);
      gj_testConfigure_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  merge  transition  place  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	73 
    -- CP-element group 288:  members (4) 
      -- CP-element group 288: 	 branch_block_stmt_33/merge_stmt_306__exit__
      -- CP-element group 288: 	 branch_block_stmt_33/assign_stmt_314_to_assign_stmt_500__entry__
      -- CP-element group 288: 	 branch_block_stmt_33/merge_stmt_306_PhiAck/$exit
      -- CP-element group 288: 	 branch_block_stmt_33/merge_stmt_306_PhiAck/phi_stmt_307_ack
      -- 
    phi_stmt_307_ack_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_307_ack_0, ack => testConfigure_CP_0_elements(288)); -- 
    -- CP-element group 289:  merge  branch  transition  place  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	120 
    -- CP-element group 289: 	166 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	122 
    -- CP-element group 289: 	123 
    -- CP-element group 289:  members (17) 
      -- CP-element group 289: 	 branch_block_stmt_33/merge_stmt_509__exit__
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_515_to_assign_stmt_521__entry__
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_515_to_assign_stmt_521__exit__
      -- CP-element group 289: 	 branch_block_stmt_33/if_stmt_522__entry__
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_515_to_assign_stmt_521/$entry
      -- CP-element group 289: 	 branch_block_stmt_33/assign_stmt_515_to_assign_stmt_521/$exit
      -- CP-element group 289: 	 branch_block_stmt_33/if_stmt_522_dead_link/$entry
      -- CP-element group 289: 	 branch_block_stmt_33/if_stmt_522_eval_test/$entry
      -- CP-element group 289: 	 branch_block_stmt_33/if_stmt_522_eval_test/$exit
      -- CP-element group 289: 	 branch_block_stmt_33/if_stmt_522_eval_test/branch_req
      -- CP-element group 289: 	 branch_block_stmt_33/R_cmp124208_523_place
      -- CP-element group 289: 	 branch_block_stmt_33/if_stmt_522_if_link/$entry
      -- CP-element group 289: 	 branch_block_stmt_33/if_stmt_522_else_link/$entry
      -- CP-element group 289: 	 branch_block_stmt_33/merge_stmt_509_PhiReqMerge
      -- CP-element group 289: 	 branch_block_stmt_33/merge_stmt_509_PhiAck/$entry
      -- CP-element group 289: 	 branch_block_stmt_33/merge_stmt_509_PhiAck/$exit
      -- CP-element group 289: 	 branch_block_stmt_33/merge_stmt_509_PhiAck/dummy
      -- 
    branch_req_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => if_stmt_522_branch_req_0); -- 
    testConfigure_CP_0_elements(289) <= OrReduce(testConfigure_CP_0_elements(120) & testConfigure_CP_0_elements(166));
    -- CP-element group 290:  transition  output  delay-element  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	125 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	294 
    -- CP-element group 290:  members (5) 
      -- CP-element group 290: 	 branch_block_stmt_33/bbx_xnph215_forx_xbody67_PhiReq/$exit
      -- CP-element group 290: 	 branch_block_stmt_33/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_564/$exit
      -- CP-element group 290: 	 branch_block_stmt_33/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/$exit
      -- CP-element group 290: 	 branch_block_stmt_33/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_568_konst_delay_trans
      -- CP-element group 290: 	 branch_block_stmt_33/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_req
      -- 
    phi_stmt_564_req_3072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_564_req_3072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(290), ack => phi_stmt_564_req_0); -- 
    -- Element group testConfigure_CP_0_elements(290) is a control-delay.
    cp_element_290_delay: control_delay_element  generic map(name => " 290_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(125), ack => testConfigure_CP_0_elements(290), clk => clk, reset =>reset);
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	167 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (2) 
      -- CP-element group 291: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/SplitProtocol/Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/SplitProtocol/Sample/ra
      -- 
    ra_3092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_570_inst_ack_0, ack => testConfigure_CP_0_elements(291)); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	167 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (2) 
      -- CP-element group 292: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/SplitProtocol/Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/SplitProtocol/Update/ca
      -- 
    ca_3097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_570_inst_ack_1, ack => testConfigure_CP_0_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/$exit
      -- CP-element group 293: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/$exit
      -- CP-element group 293: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/$exit
      -- CP-element group 293: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/$exit
      -- CP-element group 293: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_sources/type_cast_570/SplitProtocol/$exit
      -- CP-element group 293: 	 branch_block_stmt_33/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_564/phi_stmt_564_req
      -- 
    phi_stmt_564_req_3098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_564_req_3098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => phi_stmt_564_req_1); -- 
    testConfigure_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(291) & testConfigure_CP_0_elements(292);
      gj_testConfigure_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  merge  transition  place  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	290 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (2) 
      -- CP-element group 294: 	 branch_block_stmt_33/merge_stmt_563_PhiReqMerge
      -- CP-element group 294: 	 branch_block_stmt_33/merge_stmt_563_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(294) <= OrReduce(testConfigure_CP_0_elements(290) & testConfigure_CP_0_elements(293));
    -- CP-element group 295:  fork  transition  place  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	126 
    -- CP-element group 295: 	127 
    -- CP-element group 295: 	129 
    -- CP-element group 295: 	130 
    -- CP-element group 295: 	133 
    -- CP-element group 295: 	137 
    -- CP-element group 295: 	141 
    -- CP-element group 295: 	145 
    -- CP-element group 295: 	149 
    -- CP-element group 295: 	153 
    -- CP-element group 295: 	157 
    -- CP-element group 295: 	161 
    -- CP-element group 295: 	164 
    -- CP-element group 295:  members (56) 
      -- CP-element group 295: 	 branch_block_stmt_33/merge_stmt_563__exit__
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726__entry__
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_resized_1
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_scaled_1
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_computed_1
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_resize_1/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_resize_1/$exit
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_resize_1/index_resize_req
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_resize_1/index_resize_ack
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_scale_1/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_scale_1/$exit
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_scale_1/scale_rename_req
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_index_scale_1/scale_rename_ack
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_final_index_sum_regn_update_start
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_final_index_sum_regn_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_final_index_sum_regn_Sample/req
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_final_index_sum_regn_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/array_obj_ref_576_final_index_sum_regn_Update/req
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/addr_of_577_complete/req
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_sample_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/RPIPE_ConvTranspose_input_pipe_580_Sample/rr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_584_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_597_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_615_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_633_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_651_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_669_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_687_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/type_cast_705_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Update/word_access_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Update/word_access_complete/word_0/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/assign_stmt_578_to_assign_stmt_726/ptr_deref_713_Update/word_access_complete/word_0/cr
      -- CP-element group 295: 	 branch_block_stmt_33/merge_stmt_563_PhiAck/$exit
      -- CP-element group 295: 	 branch_block_stmt_33/merge_stmt_563_PhiAck/phi_stmt_564_ack
      -- 
    phi_stmt_564_ack_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_564_ack_0, ack => testConfigure_CP_0_elements(295)); -- 
    req_1635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => array_obj_ref_576_index_offset_req_0); -- 
    req_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => array_obj_ref_576_index_offset_req_1); -- 
    req_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => addr_of_577_final_reg_req_1); -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => RPIPE_ConvTranspose_input_pipe_580_inst_req_0); -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_584_inst_req_1); -- 
    cr_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_597_inst_req_1); -- 
    cr_1739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_615_inst_req_1); -- 
    cr_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_633_inst_req_1); -- 
    cr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_651_inst_req_1); -- 
    cr_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_669_inst_req_1); -- 
    cr_1851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_687_inst_req_1); -- 
    cr_1879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_705_inst_req_1); -- 
    cr_1929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => ptr_deref_713_store_0_req_1); -- 
    -- CP-element group 296:  transition  output  delay-element  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	169 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	300 
    -- CP-element group 296:  members (5) 
      -- CP-element group 296: 	 branch_block_stmt_33/bbx_xnph210_forx_xbody126_PhiReq/$exit
      -- CP-element group 296: 	 branch_block_stmt_33/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_774/$exit
      -- CP-element group 296: 	 branch_block_stmt_33/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/$exit
      -- CP-element group 296: 	 branch_block_stmt_33/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_778_konst_delay_trans
      -- CP-element group 296: 	 branch_block_stmt_33/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_req
      -- 
    phi_stmt_774_req_3126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_774_req_3126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(296), ack => phi_stmt_774_req_0); -- 
    -- Element group testConfigure_CP_0_elements(296) is a control-delay.
    cp_element_296_delay: control_delay_element  generic map(name => " 296_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(169), ack => testConfigure_CP_0_elements(296), clk => clk, reset =>reset);
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	211 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (2) 
      -- CP-element group 297: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/SplitProtocol/Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/SplitProtocol/Sample/ra
      -- 
    ra_3146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_780_inst_ack_0, ack => testConfigure_CP_0_elements(297)); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	211 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (2) 
      -- CP-element group 298: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/SplitProtocol/Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/SplitProtocol/Update/ca
      -- 
    ca_3151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_780_inst_ack_1, ack => testConfigure_CP_0_elements(298)); -- 
    -- CP-element group 299:  join  transition  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/$exit
      -- CP-element group 299: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/$exit
      -- CP-element group 299: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/$exit
      -- CP-element group 299: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/$exit
      -- CP-element group 299: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_sources/type_cast_780/SplitProtocol/$exit
      -- CP-element group 299: 	 branch_block_stmt_33/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_774/phi_stmt_774_req
      -- 
    phi_stmt_774_req_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_774_req_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(299), ack => phi_stmt_774_req_1); -- 
    testConfigure_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(297) & testConfigure_CP_0_elements(298);
      gj_testConfigure_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  merge  transition  place  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	296 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (2) 
      -- CP-element group 300: 	 branch_block_stmt_33/merge_stmt_773_PhiReqMerge
      -- CP-element group 300: 	 branch_block_stmt_33/merge_stmt_773_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(300) <= OrReduce(testConfigure_CP_0_elements(296) & testConfigure_CP_0_elements(299));
    -- CP-element group 301:  fork  transition  place  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	170 
    -- CP-element group 301: 	171 
    -- CP-element group 301: 	173 
    -- CP-element group 301: 	174 
    -- CP-element group 301: 	177 
    -- CP-element group 301: 	181 
    -- CP-element group 301: 	185 
    -- CP-element group 301: 	189 
    -- CP-element group 301: 	193 
    -- CP-element group 301: 	197 
    -- CP-element group 301: 	201 
    -- CP-element group 301: 	205 
    -- CP-element group 301: 	208 
    -- CP-element group 301:  members (56) 
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_33/merge_stmt_773__exit__
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936__entry__
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_897_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_915_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_861_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Update/word_access_complete/word_0/cr
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Update/word_access_complete/word_0/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Update/word_access_complete/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_879_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/ptr_deref_923_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_resized_1
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_scaled_1
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_computed_1
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_resize_1/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_resize_1/$exit
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_resize_1/index_resize_req
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_resize_1/index_resize_ack
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_scale_1/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_scale_1/$exit
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_scale_1/scale_rename_req
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_index_scale_1/scale_rename_ack
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_final_index_sum_regn_update_start
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_final_index_sum_regn_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_final_index_sum_regn_Sample/req
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_final_index_sum_regn_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/array_obj_ref_786_final_index_sum_regn_Update/req
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_complete/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/addr_of_787_complete/req
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/RPIPE_ConvTranspose_input_pipe_790_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_794_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_807_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_825_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_33/assign_stmt_788_to_assign_stmt_936/type_cast_843_update_start_
      -- CP-element group 301: 	 branch_block_stmt_33/merge_stmt_773_PhiAck/$exit
      -- CP-element group 301: 	 branch_block_stmt_33/merge_stmt_773_PhiAck/phi_stmt_774_ack
      -- 
    phi_stmt_774_ack_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_774_ack_0, ack => testConfigure_CP_0_elements(301)); -- 
    cr_2154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_861_inst_req_1); -- 
    cr_2210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_897_inst_req_1); -- 
    cr_2238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_915_inst_req_1); -- 
    cr_2288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => ptr_deref_923_store_0_req_1); -- 
    cr_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_879_inst_req_1); -- 
    cr_2126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_843_inst_req_1); -- 
    req_1994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => array_obj_ref_786_index_offset_req_0); -- 
    req_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => array_obj_ref_786_index_offset_req_1); -- 
    req_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => addr_of_787_final_reg_req_1); -- 
    rr_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => RPIPE_ConvTranspose_input_pipe_790_inst_req_0); -- 
    cr_2042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_794_inst_req_1); -- 
    cr_2070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_807_inst_req_1); -- 
    cr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_825_inst_req_1); -- 
    -- CP-element group 302:  merge  place  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	122 
    -- CP-element group 302: 	210 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (1) 
      -- CP-element group 302: 	 branch_block_stmt_33/merge_stmt_945_PhiReqMerge
      -- 
    testConfigure_CP_0_elements(302) <= OrReduce(testConfigure_CP_0_elements(122) & testConfigure_CP_0_elements(210));
    -- CP-element group 303:  join  fork  transition  place  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	212 
    -- CP-element group 303: 	213 
    -- CP-element group 303: 	214 
    -- CP-element group 303: 	215 
    -- CP-element group 303: 	216 
    -- CP-element group 303: 	217 
    -- CP-element group 303:  members (84) 
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_33/merge_stmt_945__exit__
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997__entry__
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_base_address_resized
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Sample/word_access_start/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_word_addrgen/root_register_ack
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Sample/word_access_start/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_update_start_
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_base_address_resized
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/word_access_complete/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Sample/word_access_start/word_0/rr
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_word_addrgen/root_register_ack
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Sample/word_access_start/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Sample/word_access_start/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Sample/word_access_start/word_0/rr
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/word_access_complete/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_update_start_
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_word_addrgen/root_register_ack
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_base_address_resized
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_update_start_
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/word_access_complete/word_0/cr
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/word_access_complete/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/word_access_complete/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/word_access_complete/word_0/cr
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_980_Update/word_access_complete/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Sample/word_access_start/word_0/rr
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Sample/word_access_start/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/word_access_complete/word_0/cr
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_956_Update/word_access_complete/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/assign_stmt_953_to_assign_stmt_997/ptr_deref_968_Sample/word_access_start/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/merge_stmt_945_PhiAck/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/merge_stmt_945_PhiAck/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/merge_stmt_945_PhiAck/dummy
      -- 
    rr_2444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_980_load_0_req_0); -- 
    rr_2344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_956_load_0_req_0); -- 
    cr_2405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_968_load_0_req_1); -- 
    cr_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_980_load_0_req_1); -- 
    rr_2394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_968_load_0_req_0); -- 
    cr_2355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_956_load_0_req_1); -- 
    testConfigure_CP_0_elements(303) <= testConfigure_CP_0_elements(302);
    -- CP-element group 304:  transition  output  delay-element  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	222 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	308 
    -- CP-element group 304:  members (5) 
      -- CP-element group 304: 	 branch_block_stmt_33/bbx_xnph_forx_xbody193_PhiReq/$exit
      -- CP-element group 304: 	 branch_block_stmt_33/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1042/$exit
      -- CP-element group 304: 	 branch_block_stmt_33/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/$exit
      -- CP-element group 304: 	 branch_block_stmt_33/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1046_konst_delay_trans
      -- CP-element group 304: 	 branch_block_stmt_33/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_req
      -- 
    phi_stmt_1042_req_3203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1042_req_3203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(304), ack => phi_stmt_1042_req_0); -- 
    -- Element group testConfigure_CP_0_elements(304) is a control-delay.
    cp_element_304_delay: control_delay_element  generic map(name => " 304_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(222), ack => testConfigure_CP_0_elements(304), clk => clk, reset =>reset);
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	231 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (2) 
      -- CP-element group 305: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/SplitProtocol/Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/SplitProtocol/Sample/ra
      -- 
    ra_3223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1048_inst_ack_0, ack => testConfigure_CP_0_elements(305)); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	231 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (2) 
      -- CP-element group 306: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/SplitProtocol/Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/SplitProtocol/Update/ca
      -- 
    ca_3228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1048_inst_ack_1, ack => testConfigure_CP_0_elements(306)); -- 
    -- CP-element group 307:  join  transition  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/$exit
      -- CP-element group 307: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/$exit
      -- CP-element group 307: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/$exit
      -- CP-element group 307: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/$exit
      -- CP-element group 307: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_sources/type_cast_1048/SplitProtocol/$exit
      -- CP-element group 307: 	 branch_block_stmt_33/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1042/phi_stmt_1042_req
      -- 
    phi_stmt_1042_req_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1042_req_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(307), ack => phi_stmt_1042_req_1); -- 
    testConfigure_cp_element_group_307: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_307"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(305) & testConfigure_CP_0_elements(306);
      gj_testConfigure_cp_element_group_307 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(307), clk => clk, reset => reset); --
    end block;
    -- CP-element group 308:  merge  transition  place  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	304 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (2) 
      -- CP-element group 308: 	 branch_block_stmt_33/merge_stmt_1041_PhiReqMerge
      -- CP-element group 308: 	 branch_block_stmt_33/merge_stmt_1041_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(308) <= OrReduce(testConfigure_CP_0_elements(304) & testConfigure_CP_0_elements(307));
    -- CP-element group 309:  fork  transition  place  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	223 
    -- CP-element group 309: 	224 
    -- CP-element group 309: 	226 
    -- CP-element group 309: 	228 
    -- CP-element group 309:  members (29) 
      -- CP-element group 309: 	 branch_block_stmt_33/merge_stmt_1041__exit__
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072__entry__
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_scale_1/scale_rename_ack
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_scale_1/scale_rename_req
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_scale_1/$exit
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_scale_1/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_resize_1/index_resize_ack
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_final_index_sum_regn_Update/req
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_resize_1/index_resize_req
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_resize_1/$exit
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_final_index_sum_regn_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_resize_1/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_computed_1
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_complete/req
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_final_index_sum_regn_Sample/req
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_final_index_sum_regn_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_scaled_1
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_final_index_sum_regn_update_start
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/array_obj_ref_1054_index_resized_1
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_complete/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_update_start_
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/addr_of_1055_update_start_
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Update/word_access_complete/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Update/word_access_complete/word_0/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/assign_stmt_1056_to_assign_stmt_1072/ptr_deref_1058_Update/word_access_complete/word_0/cr
      -- CP-element group 309: 	 branch_block_stmt_33/merge_stmt_1041_PhiAck/$exit
      -- CP-element group 309: 	 branch_block_stmt_33/merge_stmt_1041_PhiAck/phi_stmt_1042_ack
      -- 
    phi_stmt_1042_ack_3234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1042_ack_0, ack => testConfigure_CP_0_elements(309)); -- 
    req_2530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => array_obj_ref_1054_index_offset_req_1); -- 
    req_2545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => addr_of_1055_final_reg_req_1); -- 
    req_2525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => array_obj_ref_1054_index_offset_req_0); -- 
    cr_2595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => ptr_deref_1058_store_0_req_1); -- 
    -- CP-element group 310:  merge  fork  transition  place  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	220 
    -- CP-element group 310: 	230 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	232 
    -- CP-element group 310: 	233 
    -- CP-element group 310:  members (13) 
      -- CP-element group 310: 	 branch_block_stmt_33/merge_stmt_1081__exit__
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_1085__entry__
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_1085/$entry
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_update_start_
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_Sample/rr
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_33/assign_stmt_1085/type_cast_1084_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_33/merge_stmt_1081_PhiReqMerge
      -- CP-element group 310: 	 branch_block_stmt_33/merge_stmt_1081_PhiAck/$entry
      -- CP-element group 310: 	 branch_block_stmt_33/merge_stmt_1081_PhiAck/$exit
      -- CP-element group 310: 	 branch_block_stmt_33/merge_stmt_1081_PhiAck/dummy
      -- 
    rr_2626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(310), ack => type_cast_1084_inst_req_0); -- 
    cr_2631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(310), ack => type_cast_1084_inst_req_1); -- 
    testConfigure_CP_0_elements(310) <= OrReduce(testConfigure_CP_0_elements(220) & testConfigure_CP_0_elements(230));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar240_785_resized : std_logic_vector(10 downto 0);
    signal R_indvar240_785_scaled : std_logic_vector(10 downto 0);
    signal R_indvar250_575_resized : std_logic_vector(13 downto 0);
    signal R_indvar250_575_scaled : std_logic_vector(13 downto 0);
    signal R_indvar260_273_resized : std_logic_vector(0 downto 0);
    signal R_indvar260_273_scaled : std_logic_vector(0 downto 0);
    signal R_indvar263_204_resized : std_logic_vector(6 downto 0);
    signal R_indvar263_204_scaled : std_logic_vector(6 downto 0);
    signal R_indvar268_101_resized : std_logic_vector(6 downto 0);
    signal R_indvar268_101_scaled : std_logic_vector(6 downto 0);
    signal R_indvar_1053_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1053_scaled : std_logic_vector(13 downto 0);
    signal STORE_padding_312_data_0 : std_logic_vector(15 downto 0);
    signal STORE_padding_312_word_address_0 : std_logic_vector(0 downto 0);
    signal add104_693 : std_logic_vector(63 downto 0);
    signal add110_711 : std_logic_vector(63 downto 0);
    signal add136_813 : std_logic_vector(63 downto 0);
    signal add142_831 : std_logic_vector(63 downto 0);
    signal add148_849 : std_logic_vector(63 downto 0);
    signal add154_867 : std_logic_vector(63 downto 0);
    signal add160_885 : std_logic_vector(63 downto 0);
    signal add166_903 : std_logic_vector(63 downto 0);
    signal add172_921 : std_logic_vector(63 downto 0);
    signal add80_621 : std_logic_vector(63 downto 0);
    signal add86_639 : std_logic_vector(63 downto 0);
    signal add92_657 : std_logic_vector(63 downto 0);
    signal add98_675 : std_logic_vector(63 downto 0);
    signal add_603 : std_logic_vector(63 downto 0);
    signal array_obj_ref_102_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_102_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_102_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_102_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_102_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_102_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1054_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1054_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1054_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1054_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1054_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1054_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_205_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_205_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_205_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_205_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_205_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_205_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_274_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_274_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_274_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_274_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_576_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_576_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_576_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_576_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_576_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_576_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_786_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_786_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_786_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_786_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_786_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_786_root_address : std_logic_vector(10 downto 0);
    signal arrayidx114_578 : std_logic_vector(31 downto 0);
    signal arrayidx176_788 : std_logic_vector(31 downto 0);
    signal arrayidx196_1056 : std_logic_vector(31 downto 0);
    signal arrayidx19_207 : std_logic_vector(31 downto 0);
    signal arrayidx33_276 : std_logic_vector(31 downto 0);
    signal arrayidx_104 : std_logic_vector(31 downto 0);
    signal call101_684 : std_logic_vector(7 downto 0);
    signal call107_702 : std_logic_vector(7 downto 0);
    signal call129_791 : std_logic_vector(7 downto 0);
    signal call133_804 : std_logic_vector(7 downto 0);
    signal call139_822 : std_logic_vector(7 downto 0);
    signal call145_840 : std_logic_vector(7 downto 0);
    signal call151_858 : std_logic_vector(7 downto 0);
    signal call157_876 : std_logic_vector(7 downto 0);
    signal call15_210 : std_logic_vector(7 downto 0);
    signal call163_894 : std_logic_vector(7 downto 0);
    signal call169_912 : std_logic_vector(7 downto 0);
    signal call29217_251 : std_logic_vector(7 downto 0);
    signal call29_283 : std_logic_vector(7 downto 0);
    signal call3228_60 : std_logic_vector(7 downto 0);
    signal call3_132 : std_logic_vector(7 downto 0);
    signal call40_317 : std_logic_vector(7 downto 0);
    signal call42_336 : std_logic_vector(7 downto 0);
    signal call44_355 : std_logic_vector(7 downto 0);
    signal call69_581 : std_logic_vector(7 downto 0);
    signal call72_594 : std_logic_vector(7 downto 0);
    signal call77_612 : std_logic_vector(7 downto 0);
    signal call83_630 : std_logic_vector(7 downto 0);
    signal call89_648 : std_logic_vector(7 downto 0);
    signal call95_666 : std_logic_vector(7 downto 0);
    signal call_36 : std_logic_vector(7 downto 0);
    signal cmp12223_173 : std_logic_vector(0 downto 0);
    signal cmp124208_521 : std_logic_vector(0 downto 0);
    signal cmp12_239 : std_logic_vector(0 downto 0);
    signal cmp191204_997 : std_logic_vector(0 downto 0);
    signal cmp227_57 : std_logic_vector(0 downto 0);
    signal cmp65213_500 : std_logic_vector(0 downto 0);
    signal cmp_129 : std_logic_vector(0 downto 0);
    signal conv103_688 : std_logic_vector(63 downto 0);
    signal conv109_706 : std_logic_vector(63 downto 0);
    signal conv130_795 : std_logic_vector(63 downto 0);
    signal conv135_808 : std_logic_vector(63 downto 0);
    signal conv141_826 : std_logic_vector(63 downto 0);
    signal conv147_844 : std_logic_vector(63 downto 0);
    signal conv153_862 : std_logic_vector(63 downto 0);
    signal conv159_880 : std_logic_vector(63 downto 0);
    signal conv165_898 : std_logic_vector(63 downto 0);
    signal conv16_214 : std_logic_vector(31 downto 0);
    signal conv171_916 : std_logic_vector(63 downto 0);
    signal conv30218_255 : std_logic_vector(15 downto 0);
    signal conv30220_265 : std_logic_vector(15 downto 0);
    signal conv30_287 : std_logic_vector(15 downto 0);
    signal conv30x_xlcssa_307 : std_logic_vector(15 downto 0);
    signal conv41_321 : std_logic_vector(31 downto 0);
    signal conv4229_64 : std_logic_vector(31 downto 0);
    signal conv4231_81 : std_logic_vector(31 downto 0);
    signal conv43_340 : std_logic_vector(31 downto 0);
    signal conv45_359 : std_logic_vector(31 downto 0);
    signal conv4_136 : std_logic_vector(31 downto 0);
    signal conv4x_xlcssa1_144 : std_logic_vector(31 downto 0);
    signal conv4x_xlcssa_151 : std_logic_vector(31 downto 0);
    signal conv51_421 : std_logic_vector(63 downto 0);
    signal conv60_488 : std_logic_vector(63 downto 0);
    signal conv70_585 : std_logic_vector(63 downto 0);
    signal conv74_598 : std_logic_vector(63 downto 0);
    signal conv79_616 : std_logic_vector(63 downto 0);
    signal conv85_634 : std_logic_vector(63 downto 0);
    signal conv91_652 : std_logic_vector(63 downto 0);
    signal conv97_670 : std_logic_vector(63 downto 0);
    signal conv_40 : std_logic_vector(31 downto 0);
    signal exitcond10_726 : std_logic_vector(0 downto 0);
    signal exitcond19_936 : std_logic_vector(0 downto 0);
    signal exitcond20_1072 : std_logic_vector(0 downto 0);
    signal exitcond_299 : std_logic_vector(0 downto 0);
    signal iNsTr_13_120 : std_logic_vector(31 downto 0);
    signal iNsTr_1_46 : std_logic_vector(31 downto 0);
    signal iNsTr_21_230 : std_logic_vector(31 downto 0);
    signal iNsTr_26_329 : std_logic_vector(31 downto 0);
    signal iNsTr_29_348 : std_logic_vector(31 downto 0);
    signal iNsTr_32_367 : std_logic_vector(31 downto 0);
    signal iNsTr_34_379 : std_logic_vector(31 downto 0);
    signal iNsTr_35_391 : std_logic_vector(31 downto 0);
    signal iNsTr_36_403 : std_logic_vector(31 downto 0);
    signal iNsTr_37_429 : std_logic_vector(31 downto 0);
    signal iNsTr_38_441 : std_logic_vector(31 downto 0);
    signal iNsTr_39_453 : std_logic_vector(31 downto 0);
    signal iNsTr_40_465 : std_logic_vector(31 downto 0);
    signal iNsTr_45_953 : std_logic_vector(31 downto 0);
    signal iNsTr_46_965 : std_logic_vector(31 downto 0);
    signal iNsTr_47_977 : std_logic_vector(31 downto 0);
    signal iNsTr_5_163 : std_logic_vector(31 downto 0);
    signal iNsTr_60_1026 : std_logic_vector(63 downto 0);
    signal inc22_200 : std_logic_vector(31 downto 0);
    signal inc_97 : std_logic_vector(31 downto 0);
    signal indvar240_774 : std_logic_vector(63 downto 0);
    signal indvar250_564 : std_logic_vector(63 downto 0);
    signal indvar260_258 : std_logic_vector(63 downto 0);
    signal indvar263_183 : std_logic_vector(63 downto 0);
    signal indvar268_74 : std_logic_vector(63 downto 0);
    signal indvar_1042 : std_logic_vector(63 downto 0);
    signal indvarx_xnext241_931 : std_logic_vector(63 downto 0);
    signal indvarx_xnext251_721 : std_logic_vector(63 downto 0);
    signal indvarx_xnext261_293 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1067 : std_logic_vector(63 downto 0);
    signal mul184_986 : std_logic_vector(31 downto 0);
    signal mul186_991 : std_logic_vector(31 downto 0);
    signal mul50_417 : std_logic_vector(31 downto 0);
    signal mul55_474 : std_logic_vector(31 downto 0);
    signal mul57_479 : std_logic_vector(31 downto 0);
    signal mul59_484 : std_logic_vector(31 downto 0);
    signal mul_412 : std_logic_vector(31 downto 0);
    signal ptr_deref_1058_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1058_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1058_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1058_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1058_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1058_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_106_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_106_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_106_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_106_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_106_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_106_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_123_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_123_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_123_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_123_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_123_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_165_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_165_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_165_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_165_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_165_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_165_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_216_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_216_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_216_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_216_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_216_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_216_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_233_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_233_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_233_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_233_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_233_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_278_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_278_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_278_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_278_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_278_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_278_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_331_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_331_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_331_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_331_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_331_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_331_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_350_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_350_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_350_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_350_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_350_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_350_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_369_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_369_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_369_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_369_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_369_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_369_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_382_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_382_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_382_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_382_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_382_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_394_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_394_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_394_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_394_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_394_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_406_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_406_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_406_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_406_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_406_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_432_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_432_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_432_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_432_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_432_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_444_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_444_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_444_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_444_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_444_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_456_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_456_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_456_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_456_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_456_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_468_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_468_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_468_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_468_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_468_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_48_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_48_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_48_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_48_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_48_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_48_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_713_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_713_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_713_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_713_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_713_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_713_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_923_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_923_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_923_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_923_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_923_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_923_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_956_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_956_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_956_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_956_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_956_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_968_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_968_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_968_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_968_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_968_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_980_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_980_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_980_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_980_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_980_word_offset_0 : std_logic_vector(6 downto 0);
    signal shl100_681 : std_logic_vector(63 downto 0);
    signal shl106_699 : std_logic_vector(63 downto 0);
    signal shl132_801 : std_logic_vector(63 downto 0);
    signal shl138_819 : std_logic_vector(63 downto 0);
    signal shl144_837 : std_logic_vector(63 downto 0);
    signal shl150_855 : std_logic_vector(63 downto 0);
    signal shl156_873 : std_logic_vector(63 downto 0);
    signal shl162_891 : std_logic_vector(63 downto 0);
    signal shl168_909 : std_logic_vector(63 downto 0);
    signal shl76_609 : std_logic_vector(63 downto 0);
    signal shl82_627 : std_logic_vector(63 downto 0);
    signal shl88_645 : std_logic_vector(63 downto 0);
    signal shl94_663 : std_logic_vector(63 downto 0);
    signal shl_591 : std_logic_vector(63 downto 0);
    signal shr123207x_xmask_515 : std_logic_vector(63 downto 0);
    signal shr212x_xmask_494 : std_logic_vector(63 downto 0);
    signal tmp11_234 : std_logic_vector(31 downto 0);
    signal tmp12_738 : std_logic_vector(31 downto 0);
    signal tmp13_743 : std_logic_vector(31 downto 0);
    signal tmp14_748 : std_logic_vector(31 downto 0);
    signal tmp15_752 : std_logic_vector(63 downto 0);
    signal tmp16_758 : std_logic_vector(63 downto 0);
    signal tmp17_764 : std_logic_vector(0 downto 0);
    signal tmp182_957 : std_logic_vector(31 downto 0);
    signal tmp183_969 : std_logic_vector(31 downto 0);
    signal tmp185_981 : std_logic_vector(31 downto 0);
    signal tmp1_124 : std_logic_vector(31 downto 0);
    signal tmp235_1010 : std_logic_vector(31 downto 0);
    signal tmp235x_xop_1022 : std_logic_vector(31 downto 0);
    signal tmp236_1016 : std_logic_vector(0 downto 0);
    signal tmp239_1039 : std_logic_vector(63 downto 0);
    signal tmp265_224 : std_logic_vector(63 downto 0);
    signal tmp270_114 : std_logic_vector(63 downto 0);
    signal tmp3_196 : std_logic_vector(63 downto 0);
    signal tmp47_383 : std_logic_vector(31 downto 0);
    signal tmp48_395 : std_logic_vector(31 downto 0);
    signal tmp49_407 : std_logic_vector(31 downto 0);
    signal tmp53_433 : std_logic_vector(31 downto 0);
    signal tmp54_445 : std_logic_vector(31 downto 0);
    signal tmp56_457 : std_logic_vector(31 downto 0);
    signal tmp58_469 : std_logic_vector(31 downto 0);
    signal tmp5_533 : std_logic_vector(31 downto 0);
    signal tmp6_538 : std_logic_vector(31 downto 0);
    signal tmp7_542 : std_logic_vector(63 downto 0);
    signal tmp8_548 : std_logic_vector(63 downto 0);
    signal tmp9_554 : std_logic_vector(0 downto 0);
    signal tmp_93 : std_logic_vector(63 downto 0);
    signal type_cast_1008_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1014_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1020_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1030_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1037_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1046_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1048_wire : std_logic_vector(63 downto 0);
    signal type_cast_1060_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1065_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_112_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_147_wire : std_logic_vector(31 downto 0);
    signal type_cast_154_wire : std_logic_vector(31 downto 0);
    signal type_cast_156_wire : std_logic_vector(31 downto 0);
    signal type_cast_171_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_186_wire : std_logic_vector(63 downto 0);
    signal type_cast_189_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_194_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_222_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_262_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_264_wire : std_logic_vector(63 downto 0);
    signal type_cast_268_wire : std_logic_vector(15 downto 0);
    signal type_cast_270_wire : std_logic_vector(15 downto 0);
    signal type_cast_291_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_297_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_310_wire : std_logic_vector(15 downto 0);
    signal type_cast_492_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_498_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_519_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_546_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_54_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_552_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_559_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_568_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_570_wire : std_logic_vector(63 downto 0);
    signal type_cast_589_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_607_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_625_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_643_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_661_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_679_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_697_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_719_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_762_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_769_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_778_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_77_wire : std_logic_vector(63 downto 0);
    signal type_cast_780_wire : std_logic_vector(63 downto 0);
    signal type_cast_799_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_80_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_817_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_835_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_84_wire : std_logic_vector(31 downto 0);
    signal type_cast_853_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_86_wire : std_logic_vector(31 downto 0);
    signal type_cast_871_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_889_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_907_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_91_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_929_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_995_wire_constant : std_logic_vector(31 downto 0);
    signal umax18_771 : std_logic_vector(63 downto 0);
    signal umax_561 : std_logic_vector(63 downto 0);
    signal xx_xop_1032 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_padding_312_word_address_0 <= "0";
    array_obj_ref_102_constant_part_of_offset <= "0000010";
    array_obj_ref_102_offset_scale_factor_0 <= "1000000";
    array_obj_ref_102_offset_scale_factor_1 <= "0000001";
    array_obj_ref_102_resized_base_address <= "0000000";
    array_obj_ref_1054_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1054_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1054_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1054_resized_base_address <= "00000000000000";
    array_obj_ref_205_constant_part_of_offset <= "0000010";
    array_obj_ref_205_offset_scale_factor_0 <= "1000000";
    array_obj_ref_205_offset_scale_factor_1 <= "0000001";
    array_obj_ref_205_resized_base_address <= "0000000";
    array_obj_ref_274_offset_scale_factor_0 <= "1";
    array_obj_ref_274_resized_base_address <= "0";
    array_obj_ref_576_constant_part_of_offset <= "00000000000000";
    array_obj_ref_576_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_576_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_576_resized_base_address <= "00000000000000";
    array_obj_ref_786_constant_part_of_offset <= "00000100001";
    array_obj_ref_786_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_786_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_786_resized_base_address <= "00000000000";
    iNsTr_13_120 <= "00000000000000000000000000000001";
    iNsTr_1_46 <= "00000000000000000000000000000001";
    iNsTr_21_230 <= "00000000000000000000000000000001";
    iNsTr_26_329 <= "00000000000000000000000000000010";
    iNsTr_29_348 <= "00000000000000000000000000000011";
    iNsTr_32_367 <= "00000000000000000000000000000100";
    iNsTr_34_379 <= "00000000000000000000000000000010";
    iNsTr_35_391 <= "00000000000000000000000000000011";
    iNsTr_36_403 <= "00000000000000000000000000000100";
    iNsTr_37_429 <= "00000000000000000000000000000010";
    iNsTr_38_441 <= "00000000000000000000000000000011";
    iNsTr_39_453 <= "00000000000000000000000000000100";
    iNsTr_40_465 <= "00000000000000000000000000000101";
    iNsTr_45_953 <= "00000000000000000000000000000010";
    iNsTr_46_965 <= "00000000000000000000000000000011";
    iNsTr_47_977 <= "00000000000000000000000000000100";
    iNsTr_5_163 <= "00000000000000000000000000000001";
    ptr_deref_1058_word_offset_0 <= "00000000000000";
    ptr_deref_106_word_offset_0 <= "0000000";
    ptr_deref_123_word_offset_0 <= "0000000";
    ptr_deref_165_word_offset_0 <= "0000000";
    ptr_deref_216_word_offset_0 <= "0000000";
    ptr_deref_233_word_offset_0 <= "0000000";
    ptr_deref_278_word_offset_0 <= "0";
    ptr_deref_331_word_offset_0 <= "0000000";
    ptr_deref_350_word_offset_0 <= "0000000";
    ptr_deref_369_word_offset_0 <= "0000000";
    ptr_deref_382_word_offset_0 <= "0000000";
    ptr_deref_394_word_offset_0 <= "0000000";
    ptr_deref_406_word_offset_0 <= "0000000";
    ptr_deref_432_word_offset_0 <= "0000000";
    ptr_deref_444_word_offset_0 <= "0000000";
    ptr_deref_456_word_offset_0 <= "0000000";
    ptr_deref_468_word_offset_0 <= "0000000";
    ptr_deref_48_word_offset_0 <= "0000000";
    ptr_deref_713_word_offset_0 <= "00000000000000";
    ptr_deref_923_word_offset_0 <= "00000000000";
    ptr_deref_956_word_offset_0 <= "0000000";
    ptr_deref_968_word_offset_0 <= "0000000";
    ptr_deref_980_word_offset_0 <= "0000000";
    type_cast_1008_wire_constant <= "00000000000000000000000000000010";
    type_cast_1014_wire_constant <= "00000000000000000000000000000001";
    type_cast_1020_wire_constant <= "11111111111111111111111111111111";
    type_cast_1030_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1037_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1046_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1060_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1065_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_112_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_171_wire_constant <= "00000000000000000000000000000000";
    type_cast_189_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_194_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_222_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_262_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_291_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_297_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_492_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_498_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_513_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_519_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_546_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_54_wire_constant <= "00000000";
    type_cast_552_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_559_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_568_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_589_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_607_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_625_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_643_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_661_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_679_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_697_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_719_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_756_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_762_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_769_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_778_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_799_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_80_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_817_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_835_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_853_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_871_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_889_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_907_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_91_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_929_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_995_wire_constant <= "00000000000000000000000000000011";
    phi_stmt_1042: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1046_wire_constant & type_cast_1048_wire;
      req <= phi_stmt_1042_req_0 & phi_stmt_1042_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1042",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1042_ack_0,
          idata => idata,
          odata => indvar_1042,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1042
    phi_stmt_144: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_147_wire;
      req(0) <= phi_stmt_144_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_144",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_144_ack_0,
          idata => idata,
          odata => conv4x_xlcssa1_144,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_144
    phi_stmt_151: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_154_wire & type_cast_156_wire;
      req <= phi_stmt_151_req_0 & phi_stmt_151_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_151",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_151_ack_0,
          idata => idata,
          odata => conv4x_xlcssa_151,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_151
    phi_stmt_183: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_186_wire & type_cast_189_wire_constant;
      req <= phi_stmt_183_req_0 & phi_stmt_183_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_183",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_183_ack_0,
          idata => idata,
          odata => indvar263_183,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_183
    phi_stmt_258: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_262_wire_constant & type_cast_264_wire;
      req <= phi_stmt_258_req_0 & phi_stmt_258_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_258",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_258_ack_0,
          idata => idata,
          odata => indvar260_258,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_258
    phi_stmt_265: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_268_wire & type_cast_270_wire;
      req <= phi_stmt_265_req_0 & phi_stmt_265_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_265",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_265_ack_0,
          idata => idata,
          odata => conv30220_265,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_265
    phi_stmt_307: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_310_wire;
      req(0) <= phi_stmt_307_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_307",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_307_ack_0,
          idata => idata,
          odata => conv30x_xlcssa_307,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_307
    phi_stmt_564: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_568_wire_constant & type_cast_570_wire;
      req <= phi_stmt_564_req_0 & phi_stmt_564_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_564",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_564_ack_0,
          idata => idata,
          odata => indvar250_564,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_564
    phi_stmt_74: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_77_wire & type_cast_80_wire_constant;
      req <= phi_stmt_74_req_0 & phi_stmt_74_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_74",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_74_ack_0,
          idata => idata,
          odata => indvar268_74,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_74
    phi_stmt_774: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_778_wire_constant & type_cast_780_wire;
      req <= phi_stmt_774_req_0 & phi_stmt_774_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_774",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_774_ack_0,
          idata => idata,
          odata => indvar240_774,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_774
    phi_stmt_81: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_84_wire & type_cast_86_wire;
      req <= phi_stmt_81_req_0 & phi_stmt_81_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_81",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_81_ack_0,
          idata => idata,
          odata => conv4231_81,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_81
    -- flow-through select operator MUX_1038_inst
    tmp239_1039 <= xx_xop_1032 when (tmp236_1016(0) /=  '0') else type_cast_1037_wire_constant;
    -- flow-through select operator MUX_560_inst
    umax_561 <= tmp8_548 when (tmp9_554(0) /=  '0') else type_cast_559_wire_constant;
    -- flow-through select operator MUX_770_inst
    umax18_771 <= tmp16_758 when (tmp17_764(0) /=  '0') else type_cast_769_wire_constant;
    addr_of_103_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_103_final_reg_req_0;
      addr_of_103_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_103_final_reg_req_1;
      addr_of_103_final_reg_ack_1<= rack(0);
      addr_of_103_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_103_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_102_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_104,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1055_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1055_final_reg_req_0;
      addr_of_1055_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1055_final_reg_req_1;
      addr_of_1055_final_reg_ack_1<= rack(0);
      addr_of_1055_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1055_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1054_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx196_1056,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_206_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_206_final_reg_req_0;
      addr_of_206_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_206_final_reg_req_1;
      addr_of_206_final_reg_ack_1<= rack(0);
      addr_of_206_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_206_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_205_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx19_207,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_275_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_275_final_reg_req_0;
      addr_of_275_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_275_final_reg_req_1;
      addr_of_275_final_reg_ack_1<= rack(0);
      addr_of_275_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_275_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_274_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx33_276,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_577_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_577_final_reg_req_0;
      addr_of_577_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_577_final_reg_req_1;
      addr_of_577_final_reg_ack_1<= rack(0);
      addr_of_577_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_577_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_576_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx114_578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_787_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_787_final_reg_req_0;
      addr_of_787_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_787_final_reg_req_1;
      addr_of_787_final_reg_ack_1<= rack(0);
      addr_of_787_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_787_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_786_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx176_788,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1025_inst_req_0;
      type_cast_1025_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1025_inst_req_1;
      type_cast_1025_inst_ack_1<= rack(0);
      type_cast_1025_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1025_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp235x_xop_1022,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_60_1026,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1048_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1048_inst_req_0;
      type_cast_1048_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1048_inst_req_1;
      type_cast_1048_inst_ack_1<= rack(0);
      type_cast_1048_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1048_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1067,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1048_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1084_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1084_inst_req_0;
      type_cast_1084_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1084_inst_req_1;
      type_cast_1084_inst_ack_1<= rack(0);
      type_cast_1084_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1084_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul50_417,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_135_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_135_inst_req_0;
      type_cast_135_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_135_inst_req_1;
      type_cast_135_inst_ack_1<= rack(0);
      type_cast_135_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_135_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_136,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_147_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_147_inst_req_0;
      type_cast_147_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_147_inst_req_1;
      type_cast_147_inst_ack_1<= rack(0);
      type_cast_147_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_147_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_147_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_154_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_154_inst_req_0;
      type_cast_154_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_154_inst_req_1;
      type_cast_154_inst_ack_1<= rack(0);
      type_cast_154_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_154_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4229_64,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_154_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_156_inst_req_0;
      type_cast_156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_156_inst_req_1;
      type_cast_156_inst_ack_1<= rack(0);
      type_cast_156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_156_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4x_xlcssa1_144,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_156_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_186_inst_req_0;
      type_cast_186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_186_inst_req_1;
      type_cast_186_inst_ack_1<= rack(0);
      type_cast_186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp265_224,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_186_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_199_inst_req_0;
      type_cast_199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_199_inst_req_1;
      type_cast_199_inst_ack_1<= rack(0);
      type_cast_199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc22_200,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_213_inst_req_0;
      type_cast_213_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_213_inst_req_1;
      type_cast_213_inst_ack_1<= rack(0);
      type_cast_213_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_213_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_210,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_214,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_254_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_254_inst_req_0;
      type_cast_254_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_254_inst_req_1;
      type_cast_254_inst_ack_1<= rack(0);
      type_cast_254_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_254_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call29217_251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30218_255,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_264_inst_req_0;
      type_cast_264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_264_inst_req_1;
      type_cast_264_inst_ack_1<= rack(0);
      type_cast_264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_264_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext261_293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_264_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_268_inst_req_0;
      type_cast_268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_268_inst_req_1;
      type_cast_268_inst_ack_1<= rack(0);
      type_cast_268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30218_255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_268_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_270_inst_req_0;
      type_cast_270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_270_inst_req_1;
      type_cast_270_inst_ack_1<= rack(0);
      type_cast_270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_270_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30_287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_270_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_286_inst_req_0;
      type_cast_286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_286_inst_req_1;
      type_cast_286_inst_ack_1<= rack(0);
      type_cast_286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call29_283,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_310_inst_req_0;
      type_cast_310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_310_inst_req_1;
      type_cast_310_inst_ack_1<= rack(0);
      type_cast_310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30_287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_310_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_320_inst_req_0;
      type_cast_320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_320_inst_req_1;
      type_cast_320_inst_ack_1<= rack(0);
      type_cast_320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call40_317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_339_inst_req_0;
      type_cast_339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_339_inst_req_1;
      type_cast_339_inst_ack_1<= rack(0);
      type_cast_339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv43_340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_358_inst_req_0;
      type_cast_358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_358_inst_req_1;
      type_cast_358_inst_ack_1<= rack(0);
      type_cast_358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call44_355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_39_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_39_inst_req_0;
      type_cast_39_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_39_inst_req_1;
      type_cast_39_inst_ack_1<= rack(0);
      type_cast_39_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_39_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_40,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_420_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_420_inst_req_0;
      type_cast_420_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_420_inst_req_1;
      type_cast_420_inst_ack_1<= rack(0);
      type_cast_420_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_420_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul50_417,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_421,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_487_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_487_inst_req_0;
      type_cast_487_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_487_inst_req_1;
      type_cast_487_inst_ack_1<= rack(0);
      type_cast_487_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_487_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul59_484,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_488,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_541_inst_req_0;
      type_cast_541_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_541_inst_req_1;
      type_cast_541_inst_ack_1<= rack(0);
      type_cast_541_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_541_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp6_538,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp7_542,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_570_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_570_inst_req_0;
      type_cast_570_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_570_inst_req_1;
      type_cast_570_inst_ack_1<= rack(0);
      type_cast_570_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_570_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext251_721,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_570_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_584_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_584_inst_req_0;
      type_cast_584_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_584_inst_req_1;
      type_cast_584_inst_ack_1<= rack(0);
      type_cast_584_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_584_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call69_581,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_585,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_597_inst_req_0;
      type_cast_597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_597_inst_req_1;
      type_cast_597_inst_ack_1<= rack(0);
      type_cast_597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call72_594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_615_inst_req_0;
      type_cast_615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_615_inst_req_1;
      type_cast_615_inst_ack_1<= rack(0);
      type_cast_615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call77_612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_633_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_633_inst_req_0;
      type_cast_633_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_633_inst_req_1;
      type_cast_633_inst_ack_1<= rack(0);
      type_cast_633_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_633_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call83_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_634,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_63_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_63_inst_req_0;
      type_cast_63_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_63_inst_req_1;
      type_cast_63_inst_ack_1<= rack(0);
      type_cast_63_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_63_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3228_60,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4229_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_651_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_651_inst_req_0;
      type_cast_651_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_651_inst_req_1;
      type_cast_651_inst_ack_1<= rack(0);
      type_cast_651_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_651_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_652,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_669_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_669_inst_req_0;
      type_cast_669_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_669_inst_req_1;
      type_cast_669_inst_ack_1<= rack(0);
      type_cast_669_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_669_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call95_666,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv97_670,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_687_inst_req_0;
      type_cast_687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_687_inst_req_1;
      type_cast_687_inst_ack_1<= rack(0);
      type_cast_687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_688,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_705_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_705_inst_req_0;
      type_cast_705_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_705_inst_req_1;
      type_cast_705_inst_ack_1<= rack(0);
      type_cast_705_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_705_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call107_702,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_751_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_751_inst_req_0;
      type_cast_751_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_751_inst_req_1;
      type_cast_751_inst_ack_1<= rack(0);
      type_cast_751_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_751_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_77_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_77_inst_req_0;
      type_cast_77_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_77_inst_req_1;
      type_cast_77_inst_ack_1<= rack(0);
      type_cast_77_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_77_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp270_114,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_77_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_780_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_780_inst_req_0;
      type_cast_780_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_780_inst_req_1;
      type_cast_780_inst_ack_1<= rack(0);
      type_cast_780_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_780_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext241_931,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_780_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_794_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_794_inst_req_0;
      type_cast_794_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_794_inst_req_1;
      type_cast_794_inst_ack_1<= rack(0);
      type_cast_794_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_794_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_791,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_795,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_807_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_807_inst_req_0;
      type_cast_807_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_807_inst_req_1;
      type_cast_807_inst_ack_1<= rack(0);
      type_cast_807_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_807_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_804,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_808,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_825_inst_req_0;
      type_cast_825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_825_inst_req_1;
      type_cast_825_inst_ack_1<= rack(0);
      type_cast_825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call139_822,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_826,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_843_inst_req_0;
      type_cast_843_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_843_inst_req_1;
      type_cast_843_inst_ack_1<= rack(0);
      type_cast_843_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_840,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_844,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_84_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_84_inst_req_0;
      type_cast_84_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_84_inst_req_1;
      type_cast_84_inst_ack_1<= rack(0);
      type_cast_84_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_84_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_84_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_861_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_861_inst_req_0;
      type_cast_861_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_861_inst_req_1;
      type_cast_861_inst_ack_1<= rack(0);
      type_cast_861_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_861_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call151_858,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_862,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_86_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_86_inst_req_0;
      type_cast_86_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_86_inst_req_1;
      type_cast_86_inst_ack_1<= rack(0);
      type_cast_86_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_86_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4229_64,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_86_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_879_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_879_inst_req_0;
      type_cast_879_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_879_inst_req_1;
      type_cast_879_inst_ack_1<= rack(0);
      type_cast_879_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_879_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call157_876,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv159_880,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_897_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_897_inst_req_0;
      type_cast_897_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_897_inst_req_1;
      type_cast_897_inst_ack_1<= rack(0);
      type_cast_897_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_897_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call163_894,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_898,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_915_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_915_inst_req_0;
      type_cast_915_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_915_inst_req_1;
      type_cast_915_inst_ack_1<= rack(0);
      type_cast_915_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_915_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call169_912,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_916,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_96_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_96_inst_req_0;
      type_cast_96_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_96_inst_req_1;
      type_cast_96_inst_ack_1<= rack(0);
      type_cast_96_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_96_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_93,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_97,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_padding_312_gather_scatter
    process(conv30x_xlcssa_307) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv30x_xlcssa_307;
      ov(15 downto 0) := iv;
      STORE_padding_312_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_102_index_1_rename
    process(R_indvar268_101_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar268_101_resized;
      ov(6 downto 0) := iv;
      R_indvar268_101_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_102_index_1_resize
    process(indvar268_74) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar268_74;
      ov := iv(6 downto 0);
      R_indvar268_101_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_102_root_address_inst
    process(array_obj_ref_102_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_102_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_102_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1054_index_1_rename
    process(R_indvar_1053_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1053_resized;
      ov(13 downto 0) := iv;
      R_indvar_1053_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1054_index_1_resize
    process(indvar_1042) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1042;
      ov := iv(13 downto 0);
      R_indvar_1053_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1054_root_address_inst
    process(array_obj_ref_1054_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1054_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1054_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_205_index_1_rename
    process(R_indvar263_204_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar263_204_resized;
      ov(6 downto 0) := iv;
      R_indvar263_204_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_205_index_1_resize
    process(indvar263_183) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar263_183;
      ov := iv(6 downto 0);
      R_indvar263_204_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_205_root_address_inst
    process(array_obj_ref_205_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_205_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_205_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_274_index_0_rename
    process(R_indvar260_273_resized) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar260_273_resized;
      ov(0 downto 0) := iv;
      R_indvar260_273_scaled <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_274_index_0_resize
    process(indvar260_258) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar260_258;
      ov := iv(0 downto 0);
      R_indvar260_273_resized <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_274_index_offset
    process(R_indvar260_273_scaled) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar260_273_scaled;
      ov(0 downto 0) := iv;
      array_obj_ref_274_final_offset <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_274_root_address_inst
    process(array_obj_ref_274_final_offset) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_274_final_offset;
      ov(0 downto 0) := iv;
      array_obj_ref_274_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_576_index_1_rename
    process(R_indvar250_575_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar250_575_resized;
      ov(13 downto 0) := iv;
      R_indvar250_575_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_576_index_1_resize
    process(indvar250_564) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar250_564;
      ov := iv(13 downto 0);
      R_indvar250_575_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_576_root_address_inst
    process(array_obj_ref_576_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_576_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_576_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_786_index_1_rename
    process(R_indvar240_785_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar240_785_resized;
      ov(10 downto 0) := iv;
      R_indvar240_785_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_786_index_1_resize
    process(indvar240_774) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar240_774;
      ov := iv(10 downto 0);
      R_indvar240_785_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_786_root_address_inst
    process(array_obj_ref_786_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_786_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_786_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1058_addr_0
    process(ptr_deref_1058_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1058_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1058_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1058_base_resize
    process(arrayidx196_1056) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx196_1056;
      ov := iv(13 downto 0);
      ptr_deref_1058_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1058_gather_scatter
    process(type_cast_1060_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1060_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1058_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1058_root_address_inst
    process(ptr_deref_1058_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1058_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1058_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_106_addr_0
    process(ptr_deref_106_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_106_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_106_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_106_base_resize
    process(arrayidx_104) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_104;
      ov := iv(6 downto 0);
      ptr_deref_106_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_106_gather_scatter
    process(conv4231_81) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4231_81;
      ov(31 downto 0) := iv;
      ptr_deref_106_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_106_root_address_inst
    process(ptr_deref_106_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_106_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_106_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_123_addr_0
    process(ptr_deref_123_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_123_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_123_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_123_base_resize
    process(iNsTr_13_120) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_13_120;
      ov := iv(6 downto 0);
      ptr_deref_123_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_123_gather_scatter
    process(ptr_deref_123_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_123_data_0;
      ov(31 downto 0) := iv;
      tmp1_124 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_123_root_address_inst
    process(ptr_deref_123_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_123_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_123_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_165_addr_0
    process(ptr_deref_165_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_165_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_165_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_165_base_resize
    process(iNsTr_5_163) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_163;
      ov := iv(6 downto 0);
      ptr_deref_165_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_165_gather_scatter
    process(conv4x_xlcssa_151) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4x_xlcssa_151;
      ov(31 downto 0) := iv;
      ptr_deref_165_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_165_root_address_inst
    process(ptr_deref_165_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_165_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_165_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_216_addr_0
    process(ptr_deref_216_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_216_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_216_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_216_base_resize
    process(arrayidx19_207) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx19_207;
      ov := iv(6 downto 0);
      ptr_deref_216_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_216_gather_scatter
    process(conv16_214) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv16_214;
      ov(31 downto 0) := iv;
      ptr_deref_216_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_216_root_address_inst
    process(ptr_deref_216_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_216_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_216_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_233_addr_0
    process(ptr_deref_233_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_233_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_233_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_233_base_resize
    process(iNsTr_21_230) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_230;
      ov := iv(6 downto 0);
      ptr_deref_233_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_233_gather_scatter
    process(ptr_deref_233_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_233_data_0;
      ov(31 downto 0) := iv;
      tmp11_234 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_233_root_address_inst
    process(ptr_deref_233_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_233_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_233_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_addr_0
    process(ptr_deref_278_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_278_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_278_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_base_resize
    process(arrayidx33_276) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx33_276;
      ov := iv(0 downto 0);
      ptr_deref_278_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_gather_scatter
    process(conv30220_265) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv30220_265;
      ov(15 downto 0) := iv;
      ptr_deref_278_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_root_address_inst
    process(ptr_deref_278_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_278_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_278_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_331_addr_0
    process(ptr_deref_331_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_331_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_331_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_331_base_resize
    process(iNsTr_26_329) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_26_329;
      ov := iv(6 downto 0);
      ptr_deref_331_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_331_gather_scatter
    process(conv41_321) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv41_321;
      ov(31 downto 0) := iv;
      ptr_deref_331_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_331_root_address_inst
    process(ptr_deref_331_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_331_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_331_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_350_addr_0
    process(ptr_deref_350_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_350_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_350_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_350_base_resize
    process(iNsTr_29_348) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_29_348;
      ov := iv(6 downto 0);
      ptr_deref_350_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_350_gather_scatter
    process(conv43_340) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv43_340;
      ov(31 downto 0) := iv;
      ptr_deref_350_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_350_root_address_inst
    process(ptr_deref_350_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_350_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_350_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_369_addr_0
    process(ptr_deref_369_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_369_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_369_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_369_base_resize
    process(iNsTr_32_367) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_32_367;
      ov := iv(6 downto 0);
      ptr_deref_369_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_369_gather_scatter
    process(conv45_359) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv45_359;
      ov(31 downto 0) := iv;
      ptr_deref_369_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_369_root_address_inst
    process(ptr_deref_369_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_369_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_369_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_addr_0
    process(ptr_deref_382_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_382_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_382_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_base_resize
    process(iNsTr_34_379) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_34_379;
      ov := iv(6 downto 0);
      ptr_deref_382_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_gather_scatter
    process(ptr_deref_382_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_382_data_0;
      ov(31 downto 0) := iv;
      tmp47_383 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_root_address_inst
    process(ptr_deref_382_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_382_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_382_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_addr_0
    process(ptr_deref_394_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_394_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_394_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_base_resize
    process(iNsTr_35_391) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_35_391;
      ov := iv(6 downto 0);
      ptr_deref_394_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_gather_scatter
    process(ptr_deref_394_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_394_data_0;
      ov(31 downto 0) := iv;
      tmp48_395 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_root_address_inst
    process(ptr_deref_394_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_394_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_394_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_addr_0
    process(ptr_deref_406_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_406_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_base_resize
    process(iNsTr_36_403) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_36_403;
      ov := iv(6 downto 0);
      ptr_deref_406_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_gather_scatter
    process(ptr_deref_406_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_data_0;
      ov(31 downto 0) := iv;
      tmp49_407 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_root_address_inst
    process(ptr_deref_406_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_406_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_432_addr_0
    process(ptr_deref_432_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_432_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_432_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_432_base_resize
    process(iNsTr_37_429) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_429;
      ov := iv(6 downto 0);
      ptr_deref_432_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_432_gather_scatter
    process(ptr_deref_432_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_432_data_0;
      ov(31 downto 0) := iv;
      tmp53_433 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_432_root_address_inst
    process(ptr_deref_432_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_432_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_432_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_444_addr_0
    process(ptr_deref_444_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_444_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_444_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_444_base_resize
    process(iNsTr_38_441) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_38_441;
      ov := iv(6 downto 0);
      ptr_deref_444_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_444_gather_scatter
    process(ptr_deref_444_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_444_data_0;
      ov(31 downto 0) := iv;
      tmp54_445 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_444_root_address_inst
    process(ptr_deref_444_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_444_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_444_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_456_addr_0
    process(ptr_deref_456_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_456_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_456_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_456_base_resize
    process(iNsTr_39_453) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_39_453;
      ov := iv(6 downto 0);
      ptr_deref_456_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_456_gather_scatter
    process(ptr_deref_456_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_456_data_0;
      ov(31 downto 0) := iv;
      tmp56_457 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_456_root_address_inst
    process(ptr_deref_456_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_456_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_456_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_addr_0
    process(ptr_deref_468_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_468_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_468_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_base_resize
    process(iNsTr_40_465) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_40_465;
      ov := iv(6 downto 0);
      ptr_deref_468_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_gather_scatter
    process(ptr_deref_468_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_468_data_0;
      ov(31 downto 0) := iv;
      tmp58_469 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_root_address_inst
    process(ptr_deref_468_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_468_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_468_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_48_addr_0
    process(ptr_deref_48_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_48_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_48_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_48_base_resize
    process(iNsTr_1_46) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_46;
      ov := iv(6 downto 0);
      ptr_deref_48_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_48_gather_scatter
    process(conv_40) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_40;
      ov(31 downto 0) := iv;
      ptr_deref_48_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_48_root_address_inst
    process(ptr_deref_48_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_48_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_48_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_713_addr_0
    process(ptr_deref_713_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_713_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_713_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_713_base_resize
    process(arrayidx114_578) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx114_578;
      ov := iv(13 downto 0);
      ptr_deref_713_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_713_gather_scatter
    process(add110_711) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add110_711;
      ov(63 downto 0) := iv;
      ptr_deref_713_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_713_root_address_inst
    process(ptr_deref_713_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_713_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_713_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_923_addr_0
    process(ptr_deref_923_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_923_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_923_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_923_base_resize
    process(arrayidx176_788) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx176_788;
      ov := iv(10 downto 0);
      ptr_deref_923_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_923_gather_scatter
    process(add172_921) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add172_921;
      ov(63 downto 0) := iv;
      ptr_deref_923_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_923_root_address_inst
    process(ptr_deref_923_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_923_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_923_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_956_addr_0
    process(ptr_deref_956_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_956_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_956_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_956_base_resize
    process(iNsTr_45_953) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_45_953;
      ov := iv(6 downto 0);
      ptr_deref_956_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_956_gather_scatter
    process(ptr_deref_956_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_956_data_0;
      ov(31 downto 0) := iv;
      tmp182_957 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_956_root_address_inst
    process(ptr_deref_956_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_956_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_956_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_968_addr_0
    process(ptr_deref_968_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_968_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_968_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_968_base_resize
    process(iNsTr_46_965) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_46_965;
      ov := iv(6 downto 0);
      ptr_deref_968_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_968_gather_scatter
    process(ptr_deref_968_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_968_data_0;
      ov(31 downto 0) := iv;
      tmp183_969 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_968_root_address_inst
    process(ptr_deref_968_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_968_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_968_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_980_addr_0
    process(ptr_deref_980_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_980_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_980_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_980_base_resize
    process(iNsTr_47_977) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_47_977;
      ov := iv(6 downto 0);
      ptr_deref_980_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_980_gather_scatter
    process(ptr_deref_980_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_980_data_0;
      ov(31 downto 0) := iv;
      tmp185_981 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_980_root_address_inst
    process(ptr_deref_980_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_980_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_980_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1073_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond20_1072;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1073_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1073_branch_req_0,
          ack0 => if_stmt_1073_branch_ack_0,
          ack1 => if_stmt_1073_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_137_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_129;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_137_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_137_branch_req_0,
          ack0 => if_stmt_137_branch_ack_0,
          ack1 => if_stmt_137_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_174_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp12223_173;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_174_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_174_branch_req_0,
          ack0 => if_stmt_174_branch_ack_0,
          ack1 => if_stmt_174_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_240_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp12_239;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_240_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_240_branch_req_0,
          ack0 => if_stmt_240_branch_ack_0,
          ack1 => if_stmt_240_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_300_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_299;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_300_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_300_branch_req_0,
          ack0 => if_stmt_300_branch_ack_0,
          ack1 => if_stmt_300_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_501_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp65213_500;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_501_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_501_branch_req_0,
          ack0 => if_stmt_501_branch_ack_0,
          ack1 => if_stmt_501_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_522_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp124208_521;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_522_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_522_branch_req_0,
          ack0 => if_stmt_522_branch_ack_0,
          ack1 => if_stmt_522_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_65_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp227_57;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_65_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_65_branch_req_0,
          ack0 => if_stmt_65_branch_ack_0,
          ack1 => if_stmt_65_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_727_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond10_726;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_727_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_727_branch_req_0,
          ack0 => if_stmt_727_branch_ack_0,
          ack1 => if_stmt_727_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_937_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond19_936;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_937_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_937_branch_req_0,
          ack0 => if_stmt_937_branch_ack_0,
          ack1 => if_stmt_937_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_998_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp191204_997;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_998_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_998_branch_req_0,
          ack0 => if_stmt_998_branch_ack_0,
          ack1 => if_stmt_998_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1021_inst
    process(tmp235_1010) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp235_1010, type_cast_1020_wire_constant, tmp_var);
      tmp235x_xop_1022 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1031_inst
    process(iNsTr_60_1026) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_60_1026, type_cast_1030_wire_constant, tmp_var);
      xx_xop_1032 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1066_inst
    process(indvar_1042) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1042, type_cast_1065_wire_constant, tmp_var);
      indvarx_xnext_1067 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_113_inst
    process(indvar268_74) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar268_74, type_cast_112_wire_constant, tmp_var);
      tmp270_114 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_195_inst
    process(indvar263_183) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar263_183, type_cast_194_wire_constant, tmp_var);
      tmp3_196 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_223_inst
    process(indvar263_183) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar263_183, type_cast_222_wire_constant, tmp_var);
      tmp265_224 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_292_inst
    process(indvar260_258) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar260_258, type_cast_291_wire_constant, tmp_var);
      indvarx_xnext261_293 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_720_inst
    process(indvar250_564) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar250_564, type_cast_719_wire_constant, tmp_var);
      indvarx_xnext251_721 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_92_inst
    process(indvar268_74) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar268_74, type_cast_91_wire_constant, tmp_var);
      tmp_93 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_930_inst
    process(indvar240_774) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar240_774, type_cast_929_wire_constant, tmp_var);
      indvarx_xnext241_931 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_493_inst
    process(conv51_421) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv51_421, type_cast_492_wire_constant, tmp_var);
      shr212x_xmask_494 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_514_inst
    process(conv60_488) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv60_488, type_cast_513_wire_constant, tmp_var);
      shr123207x_xmask_515 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_172_inst
    process(conv4x_xlcssa_151) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv4x_xlcssa_151, type_cast_171_wire_constant, tmp_var);
      cmp12223_173 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1071_inst
    process(indvarx_xnext_1067, tmp239_1039) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1067, tmp239_1039, tmp_var);
      exitcond20_1072 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_298_inst
    process(indvarx_xnext261_293) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext261_293, type_cast_297_wire_constant, tmp_var);
      exitcond_299 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_499_inst
    process(shr212x_xmask_494) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr212x_xmask_494, type_cast_498_wire_constant, tmp_var);
      cmp65213_500 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_520_inst
    process(shr123207x_xmask_515) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr123207x_xmask_515, type_cast_519_wire_constant, tmp_var);
      cmp124208_521 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_725_inst
    process(indvarx_xnext251_721, umax_561) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext251_721, umax_561, tmp_var);
      exitcond10_726 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_935_inst
    process(indvarx_xnext241_931, umax18_771) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext241_931, umax18_771, tmp_var);
      exitcond19_936 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_55_inst
    process(call_36) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(call_36, type_cast_54_wire_constant, tmp_var);
      cmp227_57 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1009_inst
    process(mul186_991) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul186_991, type_cast_1008_wire_constant, tmp_var);
      tmp235_1010 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_547_inst
    process(tmp7_542) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp7_542, type_cast_546_wire_constant, tmp_var);
      tmp8_548 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_757_inst
    process(tmp15_752) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp15_752, type_cast_756_wire_constant, tmp_var);
      tmp16_758 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_411_inst
    process(tmp48_395, tmp47_383) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_395, tmp47_383, tmp_var);
      mul_412 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_416_inst
    process(mul_412, tmp49_407) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_412, tmp49_407, tmp_var);
      mul50_417 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_473_inst
    process(tmp54_445, tmp53_433) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_445, tmp53_433, tmp_var);
      mul55_474 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_478_inst
    process(mul55_474, tmp56_457) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul55_474, tmp56_457, tmp_var);
      mul57_479 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_483_inst
    process(mul57_479, tmp58_469) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul57_479, tmp58_469, tmp_var);
      mul59_484 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_532_inst
    process(tmp48_395, tmp47_383) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_395, tmp47_383, tmp_var);
      tmp5_533 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_537_inst
    process(tmp5_533, tmp49_407) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp5_533, tmp49_407, tmp_var);
      tmp6_538 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_737_inst
    process(tmp54_445, tmp53_433) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_445, tmp53_433, tmp_var);
      tmp12_738 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_742_inst
    process(tmp12_738, tmp56_457) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_738, tmp56_457, tmp_var);
      tmp13_743 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_747_inst
    process(tmp13_743, tmp58_469) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_743, tmp58_469, tmp_var);
      tmp14_748 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_985_inst
    process(tmp183_969, tmp182_957) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp183_969, tmp182_957, tmp_var);
      mul184_986 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_990_inst
    process(mul184_986, tmp185_981) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul184_986, tmp185_981, tmp_var);
      mul186_991 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_602_inst
    process(shl_591, conv74_598) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_591, conv74_598, tmp_var);
      add_603 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_620_inst
    process(shl76_609, conv79_616) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl76_609, conv79_616, tmp_var);
      add80_621 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_638_inst
    process(shl82_627, conv85_634) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl82_627, conv85_634, tmp_var);
      add86_639 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_656_inst
    process(shl88_645, conv91_652) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl88_645, conv91_652, tmp_var);
      add92_657 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_674_inst
    process(shl94_663, conv97_670) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl94_663, conv97_670, tmp_var);
      add98_675 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_692_inst
    process(shl100_681, conv103_688) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_681, conv103_688, tmp_var);
      add104_693 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_710_inst
    process(shl106_699, conv109_706) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl106_699, conv109_706, tmp_var);
      add110_711 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_812_inst
    process(shl132_801, conv135_808) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_801, conv135_808, tmp_var);
      add136_813 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_830_inst
    process(shl138_819, conv141_826) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl138_819, conv141_826, tmp_var);
      add142_831 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_848_inst
    process(shl144_837, conv147_844) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_837, conv147_844, tmp_var);
      add148_849 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_866_inst
    process(shl150_855, conv153_862) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl150_855, conv153_862, tmp_var);
      add154_867 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_884_inst
    process(shl156_873, conv159_880) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl156_873, conv159_880, tmp_var);
      add160_885 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_902_inst
    process(shl162_891, conv165_898) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl162_891, conv165_898, tmp_var);
      add166_903 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_920_inst
    process(shl168_909, conv171_916) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl168_909, conv171_916, tmp_var);
      add172_921 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_590_inst
    process(conv70_585) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv70_585, type_cast_589_wire_constant, tmp_var);
      shl_591 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_608_inst
    process(add_603) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_603, type_cast_607_wire_constant, tmp_var);
      shl76_609 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_626_inst
    process(add80_621) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add80_621, type_cast_625_wire_constant, tmp_var);
      shl82_627 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_644_inst
    process(add86_639) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add86_639, type_cast_643_wire_constant, tmp_var);
      shl88_645 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_662_inst
    process(add92_657) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add92_657, type_cast_661_wire_constant, tmp_var);
      shl94_663 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_680_inst
    process(add98_675) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add98_675, type_cast_679_wire_constant, tmp_var);
      shl100_681 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_698_inst
    process(add104_693) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add104_693, type_cast_697_wire_constant, tmp_var);
      shl106_699 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_800_inst
    process(conv130_795) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv130_795, type_cast_799_wire_constant, tmp_var);
      shl132_801 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_818_inst
    process(add136_813) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add136_813, type_cast_817_wire_constant, tmp_var);
      shl138_819 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_836_inst
    process(add142_831) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add142_831, type_cast_835_wire_constant, tmp_var);
      shl144_837 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_854_inst
    process(add148_849) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add148_849, type_cast_853_wire_constant, tmp_var);
      shl150_855 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_872_inst
    process(add154_867) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add154_867, type_cast_871_wire_constant, tmp_var);
      shl156_873 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_890_inst
    process(add160_885) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add160_885, type_cast_889_wire_constant, tmp_var);
      shl162_891 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_908_inst
    process(add166_903) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add166_903, type_cast_907_wire_constant, tmp_var);
      shl168_909 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1015_inst
    process(tmp235_1010) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp235_1010, type_cast_1014_wire_constant, tmp_var);
      tmp236_1016 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_996_inst
    process(mul186_991) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul186_991, type_cast_995_wire_constant, tmp_var);
      cmp191204_997 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_553_inst
    process(tmp8_548) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp8_548, type_cast_552_wire_constant, tmp_var);
      tmp9_554 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_763_inst
    process(tmp16_758) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp16_758, type_cast_762_wire_constant, tmp_var);
      tmp17_764 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_128_inst
    process(inc_97, tmp1_124) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc_97, tmp1_124, tmp_var);
      cmp_129 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_238_inst
    process(inc22_200, tmp11_234) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc22_200, tmp11_234, tmp_var);
      cmp12_239 <= tmp_var; --
    end process;
    -- shared split operator group (69) : array_obj_ref_102_index_offset 
    ApIntAdd_group_69: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar268_101_scaled;
      array_obj_ref_102_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_102_index_offset_req_0;
      array_obj_ref_102_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_102_index_offset_req_1;
      array_obj_ref_102_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_69_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_69_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_69",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000010",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : array_obj_ref_1054_index_offset 
    ApIntAdd_group_70: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1053_scaled;
      array_obj_ref_1054_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1054_index_offset_req_0;
      array_obj_ref_1054_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1054_index_offset_req_1;
      array_obj_ref_1054_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_70_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_70_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_70",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : array_obj_ref_205_index_offset 
    ApIntAdd_group_71: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar263_204_scaled;
      array_obj_ref_205_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_205_index_offset_req_0;
      array_obj_ref_205_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_205_index_offset_req_1;
      array_obj_ref_205_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_71_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_71_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_71",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000010",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : array_obj_ref_576_index_offset 
    ApIntAdd_group_72: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar250_575_scaled;
      array_obj_ref_576_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_576_index_offset_req_0;
      array_obj_ref_576_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_576_index_offset_req_1;
      array_obj_ref_576_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_72_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_72_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_72",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : array_obj_ref_786_index_offset 
    ApIntAdd_group_73: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar240_785_scaled;
      array_obj_ref_786_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_786_index_offset_req_0;
      array_obj_ref_786_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_786_index_offset_req_1;
      array_obj_ref_786_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_73_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_73_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_73",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100001",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared load operator group (0) : ptr_deref_406_load_0 ptr_deref_123_load_0 ptr_deref_382_load_0 ptr_deref_394_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_406_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_123_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_382_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_394_load_0_req_0;
      ptr_deref_406_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_123_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_382_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_394_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_406_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_123_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_382_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_394_load_0_req_1;
      ptr_deref_406_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_123_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_382_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_394_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_406_word_address_0 & ptr_deref_123_word_address_0 & ptr_deref_382_word_address_0 & ptr_deref_394_word_address_0;
      ptr_deref_406_data_0 <= data_out(127 downto 96);
      ptr_deref_123_data_0 <= data_out(95 downto 64);
      ptr_deref_382_data_0 <= data_out(63 downto 32);
      ptr_deref_394_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_456_load_0 ptr_deref_444_load_0 ptr_deref_468_load_0 ptr_deref_432_load_0 ptr_deref_233_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(34 downto 0);
      signal data_out: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2);
      -- 
    begin -- 
      reqL_unguarded(4) <= ptr_deref_456_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_444_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_468_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_432_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_233_load_0_req_0;
      ptr_deref_456_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_444_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_468_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_432_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_233_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= ptr_deref_456_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_444_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_468_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_432_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_233_load_0_req_1;
      ptr_deref_456_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_444_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_468_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_432_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_233_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_456_word_address_0 & ptr_deref_444_word_address_0 & ptr_deref_468_word_address_0 & ptr_deref_432_word_address_0 & ptr_deref_233_word_address_0;
      ptr_deref_456_data_0 <= data_out(159 downto 128);
      ptr_deref_444_data_0 <= data_out(127 downto 96);
      ptr_deref_468_data_0 <= data_out(95 downto 64);
      ptr_deref_432_data_0 <= data_out(63 downto 32);
      ptr_deref_233_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_956_load_0 ptr_deref_968_load_0 ptr_deref_980_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_956_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_968_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_980_load_0_req_0;
      ptr_deref_956_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_968_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_980_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_956_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_968_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_980_load_0_req_1;
      ptr_deref_956_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_968_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_980_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_956_word_address_0 & ptr_deref_968_word_address_0 & ptr_deref_980_word_address_0;
      ptr_deref_956_data_0 <= data_out(95 downto 64);
      ptr_deref_968_data_0 <= data_out(63 downto 32);
      ptr_deref_980_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : STORE_padding_312_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_padding_312_store_0_req_0;
      STORE_padding_312_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_padding_312_store_0_req_1;
      STORE_padding_312_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_padding_312_word_address_0;
      data_in <= STORE_padding_312_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(15 downto 0),
          mtag => memory_space_7_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1058_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1058_store_0_req_0;
      ptr_deref_1058_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1058_store_0_req_1;
      ptr_deref_1058_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1058_word_address_0;
      data_in <= ptr_deref_1058_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_48_store_0 ptr_deref_106_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_48_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_106_store_0_req_0;
      ptr_deref_48_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_106_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_48_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_106_store_0_req_1;
      ptr_deref_48_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_106_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_48_word_address_0 & ptr_deref_106_word_address_0;
      data_in <= ptr_deref_48_data_0 & ptr_deref_106_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(6 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_165_store_0 ptr_deref_216_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_165_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_216_store_0_req_0;
      ptr_deref_165_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_216_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_165_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_216_store_0_req_1;
      ptr_deref_165_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_216_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup3_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_165_word_address_0 & ptr_deref_216_word_address_0;
      data_in <= ptr_deref_165_data_0 & ptr_deref_216_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(6 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_278_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_278_store_0_req_0;
      ptr_deref_278_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_278_store_0_req_1;
      ptr_deref_278_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_278_word_address_0;
      data_in <= ptr_deref_278_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(15 downto 0),
          mtag => memory_space_8_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_331_store_0 ptr_deref_350_store_0 ptr_deref_369_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_331_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_350_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_369_store_0_req_0;
      ptr_deref_331_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_350_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_369_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_331_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_350_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_369_store_0_req_1;
      ptr_deref_331_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_350_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_369_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup5_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_331_word_address_0 & ptr_deref_350_word_address_0 & ptr_deref_369_word_address_0;
      data_in <= ptr_deref_331_data_0 & ptr_deref_350_data_0 & ptr_deref_369_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(6 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_713_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_713_store_0_req_0;
      ptr_deref_713_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_713_store_0_req_1;
      ptr_deref_713_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_713_word_address_0;
      data_in <= ptr_deref_713_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(13 downto 0),
          mdata => memory_space_4_sr_data(63 downto 0),
          mtag => memory_space_4_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_923_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_923_store_0_req_0;
      ptr_deref_923_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_923_store_0_req_1;
      ptr_deref_923_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup7_gI: SplitGuardInterface generic map(name => "StoreGroup7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_923_word_address_0;
      data_in <= ptr_deref_923_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup7 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(10 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup7 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_611_inst RPIPE_ConvTranspose_input_pipe_593_inst RPIPE_ConvTranspose_input_pipe_580_inst RPIPE_ConvTranspose_input_pipe_911_inst RPIPE_ConvTranspose_input_pipe_629_inst RPIPE_ConvTranspose_input_pipe_821_inst RPIPE_ConvTranspose_input_pipe_647_inst RPIPE_ConvTranspose_input_pipe_839_inst RPIPE_ConvTranspose_input_pipe_665_inst RPIPE_ConvTranspose_input_pipe_857_inst RPIPE_ConvTranspose_input_pipe_790_inst RPIPE_ConvTranspose_input_pipe_683_inst RPIPE_ConvTranspose_input_pipe_875_inst RPIPE_ConvTranspose_input_pipe_701_inst RPIPE_ConvTranspose_input_pipe_803_inst RPIPE_ConvTranspose_input_pipe_893_inst RPIPE_ConvTranspose_input_pipe_35_inst RPIPE_ConvTranspose_input_pipe_59_inst RPIPE_ConvTranspose_input_pipe_131_inst RPIPE_ConvTranspose_input_pipe_209_inst RPIPE_ConvTranspose_input_pipe_250_inst RPIPE_ConvTranspose_input_pipe_282_inst RPIPE_ConvTranspose_input_pipe_316_inst RPIPE_ConvTranspose_input_pipe_335_inst RPIPE_ConvTranspose_input_pipe_354_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(199 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 24 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 24 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 24 downto 0);
      signal guard_vector : std_logic_vector( 24 downto 0);
      constant outBUFs : IntegerArray(24 downto 0) := (24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(24 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false);
      constant guardBuffering: IntegerArray(24 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2);
      -- 
    begin -- 
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_611_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_593_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_580_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_911_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_629_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_821_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_647_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_839_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_665_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_857_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_790_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_683_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_875_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_701_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_803_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_893_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_131_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_209_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_250_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_282_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_335_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_354_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_611_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_593_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_580_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_911_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_629_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_821_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_647_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_839_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_665_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_857_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_790_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_683_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_875_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_701_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_803_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_893_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_131_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_209_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_250_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_282_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_335_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_354_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_611_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_593_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_580_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_911_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_629_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_821_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_647_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_839_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_665_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_857_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_790_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_683_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_875_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_701_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_803_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_893_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_131_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_209_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_250_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_282_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_335_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_354_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_611_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_593_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_580_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_911_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_629_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_821_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_647_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_839_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_665_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_857_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_790_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_683_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_875_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_701_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_803_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_893_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_131_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_209_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_250_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_282_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_335_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_354_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      call77_612 <= data_out(199 downto 192);
      call72_594 <= data_out(191 downto 184);
      call69_581 <= data_out(183 downto 176);
      call169_912 <= data_out(175 downto 168);
      call83_630 <= data_out(167 downto 160);
      call139_822 <= data_out(159 downto 152);
      call89_648 <= data_out(151 downto 144);
      call145_840 <= data_out(143 downto 136);
      call95_666 <= data_out(135 downto 128);
      call151_858 <= data_out(127 downto 120);
      call129_791 <= data_out(119 downto 112);
      call101_684 <= data_out(111 downto 104);
      call157_876 <= data_out(103 downto 96);
      call107_702 <= data_out(95 downto 88);
      call133_804 <= data_out(87 downto 80);
      call163_894 <= data_out(79 downto 72);
      call_36 <= data_out(71 downto 64);
      call3228_60 <= data_out(63 downto 56);
      call3_132 <= data_out(55 downto 48);
      call15_210 <= data_out(47 downto 40);
      call29217_251 <= data_out(39 downto 32);
      call29_283 <= data_out(31 downto 24);
      call40_317 <= data_out(23 downto 16);
      call42_336 <= data_out(15 downto 8);
      call44_355 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 25, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 25,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(5 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(5 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(41 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(119 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(5 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(5 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(191 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(11 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(79 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 21),
      memory_space_1_lr_tag => memory_space_1_lr_tag(83 downto 63),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 96),
      memory_space_1_lc_tag => memory_space_1_lc_tag(11 downto 9),
      memory_space_2_lr_req => memory_space_2_lr_req(3 downto 3),
      memory_space_2_lr_ack => memory_space_2_lr_ack(3 downto 3),
      memory_space_2_lr_addr => memory_space_2_lr_addr(27 downto 21),
      memory_space_2_lr_tag => memory_space_2_lr_tag(83 downto 63),
      memory_space_2_lc_req => memory_space_2_lc_req(3 downto 3),
      memory_space_2_lc_ack => memory_space_2_lc_ack(3 downto 3),
      memory_space_2_lc_data => memory_space_2_lc_data(127 downto 96),
      memory_space_2_lc_tag => memory_space_2_lc_tag(11 downto 9),
      memory_space_3_lr_req => memory_space_3_lr_req(3 downto 3),
      memory_space_3_lr_ack => memory_space_3_lr_ack(3 downto 3),
      memory_space_3_lr_addr => memory_space_3_lr_addr(27 downto 21),
      memory_space_3_lr_tag => memory_space_3_lr_tag(79 downto 60),
      memory_space_3_lc_req => memory_space_3_lc_req(3 downto 3),
      memory_space_3_lc_ack => memory_space_3_lc_ack(3 downto 3),
      memory_space_3_lc_data => memory_space_3_lc_data(127 downto 96),
      memory_space_3_lc_tag => memory_space_3_lc_tag(7 downto 6),
      memory_space_4_lr_req => memory_space_4_lr_req(3 downto 3),
      memory_space_4_lr_ack => memory_space_4_lr_ack(3 downto 3),
      memory_space_4_lr_addr => memory_space_4_lr_addr(55 downto 42),
      memory_space_4_lr_tag => memory_space_4_lr_tag(75 downto 57),
      memory_space_4_lc_req => memory_space_4_lc_req(3 downto 3),
      memory_space_4_lc_ack => memory_space_4_lc_ack(3 downto 3),
      memory_space_4_lc_data => memory_space_4_lc_data(255 downto 192),
      memory_space_4_lc_tag => memory_space_4_lc_tag(3 downto 3),
      memory_space_7_lr_req => memory_space_7_lr_req(3 downto 3),
      memory_space_7_lr_ack => memory_space_7_lr_ack(3 downto 3),
      memory_space_7_lr_addr => memory_space_7_lr_addr(3 downto 3),
      memory_space_7_lr_tag => memory_space_7_lr_tag(75 downto 57),
      memory_space_7_lc_req => memory_space_7_lc_req(3 downto 3),
      memory_space_7_lc_ack => memory_space_7_lc_ack(3 downto 3),
      memory_space_7_lc_data => memory_space_7_lc_data(63 downto 48),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 3),
      memory_space_8_lr_req => memory_space_8_lr_req(3 downto 3),
      memory_space_8_lr_ack => memory_space_8_lr_ack(3 downto 3),
      memory_space_8_lr_addr => memory_space_8_lr_addr(3 downto 3),
      memory_space_8_lr_tag => memory_space_8_lr_tag(79 downto 60),
      memory_space_8_lc_req => memory_space_8_lc_req(3 downto 3),
      memory_space_8_lc_ack => memory_space_8_lc_ack(3 downto 3),
      memory_space_8_lc_data => memory_space_8_lc_data(63 downto 48),
      memory_space_8_lc_tag => memory_space_8_lc_tag(7 downto 6),
      memory_space_6_sr_req => memory_space_6_sr_req(3 downto 3),
      memory_space_6_sr_ack => memory_space_6_sr_ack(3 downto 3),
      memory_space_6_sr_addr => memory_space_6_sr_addr(55 downto 42),
      memory_space_6_sr_data => memory_space_6_sr_data(255 downto 192),
      memory_space_6_sr_tag => memory_space_6_sr_tag(75 downto 57),
      memory_space_6_sc_req => memory_space_6_sc_req(3 downto 3),
      memory_space_6_sc_ack => memory_space_6_sc_ack(3 downto 3),
      memory_space_6_sc_tag => memory_space_6_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(20 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(62 downto 42),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(95 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(8 downto 6),
      memory_space_2_lr_req => memory_space_2_lr_req(2 downto 2),
      memory_space_2_lr_ack => memory_space_2_lr_ack(2 downto 2),
      memory_space_2_lr_addr => memory_space_2_lr_addr(20 downto 14),
      memory_space_2_lr_tag => memory_space_2_lr_tag(62 downto 42),
      memory_space_2_lc_req => memory_space_2_lc_req(2 downto 2),
      memory_space_2_lc_ack => memory_space_2_lc_ack(2 downto 2),
      memory_space_2_lc_data => memory_space_2_lc_data(95 downto 64),
      memory_space_2_lc_tag => memory_space_2_lc_tag(8 downto 6),
      memory_space_3_lr_req => memory_space_3_lr_req(2 downto 2),
      memory_space_3_lr_ack => memory_space_3_lr_ack(2 downto 2),
      memory_space_3_lr_addr => memory_space_3_lr_addr(20 downto 14),
      memory_space_3_lr_tag => memory_space_3_lr_tag(59 downto 40),
      memory_space_3_lc_req => memory_space_3_lc_req(2 downto 2),
      memory_space_3_lc_ack => memory_space_3_lc_ack(2 downto 2),
      memory_space_3_lc_data => memory_space_3_lc_data(95 downto 64),
      memory_space_3_lc_tag => memory_space_3_lc_tag(5 downto 4),
      memory_space_4_lr_req => memory_space_4_lr_req(2 downto 2),
      memory_space_4_lr_ack => memory_space_4_lr_ack(2 downto 2),
      memory_space_4_lr_addr => memory_space_4_lr_addr(41 downto 28),
      memory_space_4_lr_tag => memory_space_4_lr_tag(56 downto 38),
      memory_space_4_lc_req => memory_space_4_lc_req(2 downto 2),
      memory_space_4_lc_ack => memory_space_4_lc_ack(2 downto 2),
      memory_space_4_lc_data => memory_space_4_lc_data(191 downto 128),
      memory_space_4_lc_tag => memory_space_4_lc_tag(2 downto 2),
      memory_space_7_lr_req => memory_space_7_lr_req(2 downto 2),
      memory_space_7_lr_ack => memory_space_7_lr_ack(2 downto 2),
      memory_space_7_lr_addr => memory_space_7_lr_addr(2 downto 2),
      memory_space_7_lr_tag => memory_space_7_lr_tag(56 downto 38),
      memory_space_7_lc_req => memory_space_7_lc_req(2 downto 2),
      memory_space_7_lc_ack => memory_space_7_lc_ack(2 downto 2),
      memory_space_7_lc_data => memory_space_7_lc_data(47 downto 32),
      memory_space_7_lc_tag => memory_space_7_lc_tag(2 downto 2),
      memory_space_8_lr_req => memory_space_8_lr_req(2 downto 2),
      memory_space_8_lr_ack => memory_space_8_lr_ack(2 downto 2),
      memory_space_8_lr_addr => memory_space_8_lr_addr(2 downto 2),
      memory_space_8_lr_tag => memory_space_8_lr_tag(59 downto 40),
      memory_space_8_lc_req => memory_space_8_lc_req(2 downto 2),
      memory_space_8_lc_ack => memory_space_8_lc_ack(2 downto 2),
      memory_space_8_lc_data => memory_space_8_lc_data(47 downto 32),
      memory_space_8_lc_tag => memory_space_8_lc_tag(5 downto 4),
      memory_space_6_sr_req => memory_space_6_sr_req(2 downto 2),
      memory_space_6_sr_ack => memory_space_6_sr_ack(2 downto 2),
      memory_space_6_sr_addr => memory_space_6_sr_addr(41 downto 28),
      memory_space_6_sr_data => memory_space_6_sr_data(191 downto 128),
      memory_space_6_sr_tag => memory_space_6_sr_tag(56 downto 38),
      memory_space_6_sc_req => memory_space_6_sc_req(2 downto 2),
      memory_space_6_sc_ack => memory_space_6_sc_ack(2 downto 2),
      memory_space_6_sc_tag => memory_space_6_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 7),
      memory_space_1_lr_tag => memory_space_1_lr_tag(41 downto 21),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 3),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 7),
      memory_space_2_lr_tag => memory_space_2_lr_tag(41 downto 21),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(5 downto 3),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 7),
      memory_space_3_lr_tag => memory_space_3_lr_tag(39 downto 20),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 32),
      memory_space_3_lc_tag => memory_space_3_lc_tag(3 downto 2),
      memory_space_4_lr_req => memory_space_4_lr_req(1 downto 1),
      memory_space_4_lr_ack => memory_space_4_lr_ack(1 downto 1),
      memory_space_4_lr_addr => memory_space_4_lr_addr(27 downto 14),
      memory_space_4_lr_tag => memory_space_4_lr_tag(37 downto 19),
      memory_space_4_lc_req => memory_space_4_lc_req(1 downto 1),
      memory_space_4_lc_ack => memory_space_4_lc_ack(1 downto 1),
      memory_space_4_lc_data => memory_space_4_lc_data(127 downto 64),
      memory_space_4_lc_tag => memory_space_4_lc_tag(1 downto 1),
      memory_space_7_lr_req => memory_space_7_lr_req(1 downto 1),
      memory_space_7_lr_ack => memory_space_7_lr_ack(1 downto 1),
      memory_space_7_lr_addr => memory_space_7_lr_addr(1 downto 1),
      memory_space_7_lr_tag => memory_space_7_lr_tag(37 downto 19),
      memory_space_7_lc_req => memory_space_7_lc_req(1 downto 1),
      memory_space_7_lc_ack => memory_space_7_lc_ack(1 downto 1),
      memory_space_7_lc_data => memory_space_7_lc_data(31 downto 16),
      memory_space_7_lc_tag => memory_space_7_lc_tag(1 downto 1),
      memory_space_8_lr_req => memory_space_8_lr_req(1 downto 1),
      memory_space_8_lr_ack => memory_space_8_lr_ack(1 downto 1),
      memory_space_8_lr_addr => memory_space_8_lr_addr(1 downto 1),
      memory_space_8_lr_tag => memory_space_8_lr_tag(39 downto 20),
      memory_space_8_lc_req => memory_space_8_lc_req(1 downto 1),
      memory_space_8_lc_ack => memory_space_8_lc_ack(1 downto 1),
      memory_space_8_lc_data => memory_space_8_lc_data(31 downto 16),
      memory_space_8_lc_tag => memory_space_8_lc_tag(3 downto 2),
      memory_space_6_sr_req => memory_space_6_sr_req(1 downto 1),
      memory_space_6_sr_ack => memory_space_6_sr_ack(1 downto 1),
      memory_space_6_sr_addr => memory_space_6_sr_addr(27 downto 14),
      memory_space_6_sr_data => memory_space_6_sr_data(127 downto 64),
      memory_space_6_sr_tag => memory_space_6_sr_tag(37 downto 19),
      memory_space_6_sc_req => memory_space_6_sc_req(1 downto 1),
      memory_space_6_sc_ack => memory_space_6_sc_ack(1 downto 1),
      memory_space_6_sc_tag => memory_space_6_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(6 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(6 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(20 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(2 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(6 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(19 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(1 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(13 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(18 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(63 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(0 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(18 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(0 downto 0),
      memory_space_8_lr_req => memory_space_8_lr_req(0 downto 0),
      memory_space_8_lr_ack => memory_space_8_lr_ack(0 downto 0),
      memory_space_8_lr_addr => memory_space_8_lr_addr(0 downto 0),
      memory_space_8_lr_tag => memory_space_8_lr_tag(19 downto 0),
      memory_space_8_lc_req => memory_space_8_lc_req(0 downto 0),
      memory_space_8_lc_ack => memory_space_8_lc_ack(0 downto 0),
      memory_space_8_lc_data => memory_space_8_lc_data(15 downto 0),
      memory_space_8_lc_tag => memory_space_8_lc_tag(1 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(13 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(63 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(18 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(4 downto 4),
      memory_space_3_lr_ack => memory_space_3_lr_ack(4 downto 4),
      memory_space_3_lr_addr => memory_space_3_lr_addr(34 downto 28),
      memory_space_3_lr_tag => memory_space_3_lr_tag(99 downto 80),
      memory_space_3_lc_req => memory_space_3_lc_req(4 downto 4),
      memory_space_3_lc_ack => memory_space_3_lc_ack(4 downto 4),
      memory_space_3_lc_data => memory_space_3_lc_data(159 downto 128),
      memory_space_3_lc_tag => memory_space_3_lc_tag(9 downto 8),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(13 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(18 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(4 downto 4),
      memory_space_1_lr_ack => memory_space_1_lr_ack(4 downto 4),
      memory_space_1_lr_addr => memory_space_1_lr_addr(34 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(104 downto 84),
      memory_space_1_lc_req => memory_space_1_lc_req(4 downto 4),
      memory_space_1_lc_ack => memory_space_1_lc_ack(4 downto 4),
      memory_space_1_lc_data => memory_space_1_lc_data(159 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(14 downto 12),
      memory_space_2_lr_req => memory_space_2_lr_req(4 downto 4),
      memory_space_2_lr_ack => memory_space_2_lr_ack(4 downto 4),
      memory_space_2_lr_addr => memory_space_2_lr_addr(34 downto 28),
      memory_space_2_lr_tag => memory_space_2_lr_tag(104 downto 84),
      memory_space_2_lc_req => memory_space_2_lc_req(4 downto 4),
      memory_space_2_lc_ack => memory_space_2_lc_ack(4 downto 4),
      memory_space_2_lc_data => memory_space_2_lc_data(159 downto 128),
      memory_space_2_lc_tag => memory_space_2_lc_tag(14 downto 12),
      memory_space_3_lr_req => memory_space_3_lr_req(5 downto 5),
      memory_space_3_lr_ack => memory_space_3_lr_ack(5 downto 5),
      memory_space_3_lr_addr => memory_space_3_lr_addr(41 downto 35),
      memory_space_3_lr_tag => memory_space_3_lr_tag(119 downto 100),
      memory_space_3_lc_req => memory_space_3_lc_req(5 downto 5),
      memory_space_3_lc_ack => memory_space_3_lc_ack(5 downto 5),
      memory_space_3_lc_data => memory_space_3_lc_data(191 downto 160),
      memory_space_3_lc_tag => memory_space_3_lc_tag(11 downto 10),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(6 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(6 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(20 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(6 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(31 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(19 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(13 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(63 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(18 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(10 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(63 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(0 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(4 downto 4),
      memory_space_6_sr_ack => memory_space_6_sr_ack(4 downto 4),
      memory_space_6_sr_addr => memory_space_6_sr_addr(69 downto 56),
      memory_space_6_sr_data => memory_space_6_sr_data(319 downto 256),
      memory_space_6_sr_tag => memory_space_6_sr_tag(94 downto 76),
      memory_space_6_sc_req => memory_space_6_sc_req(4 downto 4),
      memory_space_6_sc_ack => memory_space_6_sc_ack(4 downto 4),
      memory_space_6_sc_tag => memory_space_6_sc_tag(4 downto 4),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(15 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(18 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(0 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(0 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(15 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(19 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 6,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_5: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
